// IWLS benchmark module "C3540.iscas" printed on Wed May 29 16:28:04 2002
module test3 (\1(0) , \13(1) , \20(2) , \33(3) , \41(4) , \45(5) , \50(6) , \58(7) , \68(8) , \77(9) , \87(10) , \97(11) , \107(12) , \116(13) , \124(14) , \125(15) , \128(16) , \132(17) , \137(18) , \143(19) , \150(20) , \159(21) , \169(22) , \179(23) , \190(24) , \200(25) , \213(26) , \222(27) , \223(28) , \226(29) , \232(30) , \238(31) , \244(32) , \250(33) , \257(34) , \264(35) , \270(36) , \274(37) , \283(38) , \294(39) , \303(40) , \311(41) , \317(42) , \322(43) , \326(44) , \329(45) , \330(46) , \343(47) , \1698(48) , \2897(49) , \353(405) , \355(399) , \361(940) , \358(1161) , \351(1247) , \372(1243) , \369(1321) , \399(1428) , \364(1484) , \396(1504) , \384(1553) , \367(1585) , \387(1616) , \393(1605) , \390(1603) , \378(1597) , \375(1624) , \381(1626) , \407(1657) , \409(1670) , \405(1717) , \402(1718) );
input
  \244(32) ,
  \50(6) ,
  \322(43) ,
  \33(3) ,
  \116(13) ,
  \326(44) ,
  \222(27) ,
  \250(33) ,
  \226(29) ,
  \58(7) ,
  \107(12) ,
  \317(42) ,
  \77(9) ,
  \213(26) ,
  \200(25) ,
  \20(2) ,
  \150(20) ,
  \41(4) ,
  \232(30) ,
  \45(5) ,
  \1698(48) ,
  \264(35) ,
  \223(28) ,
  \132(17) ,
  \68(8) ,
  \283(38) ,
  \13(1) ,
  \270(36) ,
  \274(37) ,
  \311(41) ,
  \159(21) ,
  \343(47) ,
  \1(0) ,
  \137(18) ,
  \330(46) ,
  \87(10) ,
  \124(14) ,
  \128(16) ,
  \169(22) ,
  \2897(49) ,
  \143(19) ,
  \329(45) ,
  \238(31) ,
  \97(11) ,
  \294(39) ,
  \303(40) ,
  \179(23) ,
  \190(24) ,
  \257(34) ,
  \125(15) ;
output
  \387(1616) ,
  \390(1603) ,
  \409(1670) ,
  \369(1321) ,
  \402(1718) ,
  \353(405) ,
  \375(1624) ,
  \384(1553) ,
  \407(1657) ,
  \361(940) ,
  \372(1243) ,
  \355(399) ,
  \378(1597) ,
  \393(1605) ,
  \399(1428) ,
  \364(1484) ,
  \351(1247) ,
  \358(1161) ,
  \396(1504) ,
  \405(1717) ,
  \381(1626) ,
  \367(1585) ;
wire
  \703(1187) ,
  \2580(1425) ,
  \920(361) ,
  \2886(1658) ,
  \2742(1390) ,
  \2997(1038) ,
  \574(585) ,
  \1539(1079) ,
  \2907(1683) ,
  \1476(757) ,
  \699(430) ,
  \3261(1438) ,
  \912(250) ,
  \1678(1254) ,
  \3196(1198) ,
  \2325(1204) ,
  \1940(1103) ,
  \2782(1581) ,
  \3473(1604) ,
  \3268(1414) ,
  \2654(1337) ,
  \776(107) ,
  \1677(1324) ,
  \2659(1568) ,
  \463(88) ,
  \1135(518) ,
  \784(191) ,
  \2730(1600) ,
  \1733(389) ,
  \2903(349) ,
  \2467(1275) ,
  \910(527) ,
  \1492(756) ,
  \1594(1026) ,
  \2722(1586) ,
  \2991(973) ,
  \2162(341) ,
  \1144(372) ,
  \1737(297) ,
  \985(378) ,
  \2100(1057) ,
  \1725(286) ,
  \2947(56) ,
  \1325(662) ,
  \1009(318) ,
  \1270(823) ,
  \2336(1295) ,
  \2828(1640) ,
  \896(176) ,
  \1311(613) ,
  \3411(1403) ,
  \648(526) ,
  \2669(1563) ,
  \2549(1559) ,
  \2274(1214) ,
  \1004(252) ,
  \650(273) ,
  \504(76) ,
  \927(347) ,
  \1462(686) ,
  \1385(898) ,
  \2196(1007) ,
  \[0] ,
  \2488(503) ,
  \2965(218) ,
  \2717(557) ,
  \2149(1104) ,
  \[1] ,
  \3515(1635) ,
  \[2] ,
  \2140(926) ,
  \1644(1354) ,
  \1654(582) ,
  \1652(1090) ,
  \2745(1521) ,
  \[3] ,
  \1245(705) ,
  \2214(342) ,
  \626(158) ,
  \2777(1445) ,
  \[4] ,
  \1753(290) ,
  \2163(456) ,
  \1352(865) ,
  \[5] ,
  \3017(169) ,
  \3294(1347) ,
  \[6] ,
  \613(423) ,
  \[7] ,
  \1337(895) ,
  \2337(1265) ,
  \2946(140) ,
  \[8] ,
  \1332(646) ,
  \383(1541) ,
  \[9] ,
  \3187(1176) ,
  \1266(901) ,
  \2799(1583) ,
  \955(1536) ,
  \1903(1034) ,
  \467(87) ,
  \2770(573) ,
  \2709(1587) ,
  \1494(912) ,
  \1254(831) ,
  \3197(1177) ,
  \1717(183) ,
  \3015(270) ,
  \646(248) ,
  \2058(454) ,
  \1866(900) ,
  \1306(821) ,
  \1330(710) ,
  \732(117) ,
  \3425(130) ,
  \2120(1069) ,
  \1533(421) ,
  \2934(59) ,
  \999(415) ,
  \2260(1054) ,
  \1241(673) ,
  \3345(1535) ,
  \3555(1646) ,
  \1921(495) ,
  \2380(1148) ,
  \368(1296) ,
  \984(408) ,
  \1297(628) ,
  \683(434) ,
  \1699(105) ,
  \1309(677) ,
  \2855(1679) ,
  \2883(1595) ,
  \2643(1328) ,
  \1436(870) ,
  \1657(1132) ,
  \3505(1555) ,
  \2785(468) ,
  \1333(814) ,
  \2508(1381) ,
  \3087(90) ,
  \1499(704) ,
  \1912(1076) ,
  \3353(1456) ,
  \1729(501) ,
  \2383(943) ,
  \975(321) ,
  \403(1713) ,
  \828(93) ,
  \2394(1228) ,
  \1321(802) ,
  \2057(339) ,
  \2215(457) ,
  \2982(590) ,
  \3363(1458) ,
  \3347(1434) ,
  \3153(1269) ,
  \2109(340) ,
  \3321(1406) ,
  \3371(1405) ,
  \1946(1146) ,
  \3311(1408) ,
  \2094(1002) ,
  \926(563) ,
  \2311(1109) ,
  \3228(1040) ,
  \1265(832) ,
  \618(1017) ,
  \2367(947) ,
  \1293(596) ,
  \3237(1171) ,
  \406(1643) ,
  \2930(1649) ,
  \2814(1467) ,
  \3544(1609) ,
  \2034(1009) ,
  \1336(885) ,
  \3540(1706) ,
  \2406(1284) ,
  \621(170) ,
  \3062(721) ,
  \3098(153) ,
  \1503(749) ,
  \3101(160) ,
  \1773(345) ,
  \1481(623) ,
  \1495(672) ,
  \1404(868) ,
  \1507(759) ,
  \816(179) ,
  \2257(1053) ,
  \694(435) ,
  \2906(1677) ,
  \2791(1573) ,
  \3178(1046) ,
  \3377(1433) ,
  \2863(1707) ,
  \1168(513) ,
  \2594(1526) ,
  \2661(1561) ,
  \549(139) ,
  \1313(709) ,
  \798(102) ,
  \1420(869) ,
  \1099(504) ,
  \2657(1368) ,
  \3177(1216) ,
  \692(1157) ,
  \2642(1304) ,
  \2328(1101) ,
  \630(246) ,
  \675(178) ,
  \1992(966) ,
  \1640(1289) ,
  \1978(933) ,
  \1401(776) ,
  \2698(556) ,
  \1608(1089) ,
  \691(524) ,
  \1012(386) ,
  \3044(245) ,
  \1365(632) ,
  \2975(498) ,
  \647(391) ,
  \3251(1208) ,
  \3417(1431) ,
  \3312(1290) ,
  \3093(171) ,
  \2051(104) ,
  \2046(1060) ,
  \3260(1436) ,
  \1809(343) ,
  \1716(294) ,
  \3313(1336) ,
  \1287(817) ,
  \2616(1421) ,
  \1743(496) ,
  \2324(1202) ,
  \1328(614) ,
  \2990(481) ,
  \2674(1549) ,
  \2323(1238) ,
  \1406(849) ,
  \2314(1205) ,
  \1953(452) ,
  \2273(1218) ,
  \2671(1550) ,
  \365(1570) ,
  \1628(448) ,
  \2856(1690) ,
  \3303(1340) ,
  \1808(195) ,
  \2895(1659) ,
  \2955(222) ,
  \2513(1343) ,
  \1480(607) ,
  \1589(306) ,
  \575(586) ,
  \1952(337) ,
  \1479(687) ,
  \1302(903) ,
  \3137(1222) ,
  \2887(1647) ,
  \905(155) ,
  \3435(1528) ,
  \2312(1175) ,
  \2532(1303) ,
  \1920(281) ,
  \1563(329) ,
  \1369(856) ,
  \1274(659) ,
  \2811(1393) ,
  \3127(1221) ,
  \1583(1021) ,
  \1655(437) ,
  \1873(741) ,
  \3227(1210) ,
  \2690(1611) ,
  \2706(1444) ,
  \359(587) ,
  \1281(643) ,
  \1493(753) ,
  \1588(1084) ,
  \914(440) ,
  \600(1012) ,
  \2664(1544) ,
  \2787(574) ,
  \1667(1280) ,
  \3467(1591) ,
  \2110(455) ,
  \2396(1253) ,
  \3539(1692) ,
  \587(54) ,
  \3323(1138) ,
  \1349(647) ,
  \1485(655) ,
  \3514(1634) ,
  \2432(1189) ,
  \1761(352) ,
  \1625(732) ,
  \1653(1357) ,
  \1260(610) ,
  \2957(53) ,
  \1380(697) ,
  \3045(383) ,
  \2048(1111) ,
  \2184(747) ,
  \2687(1388) ,
  \1963(881) ,
  \1347(711) ,
  \3146(1167) ,
  \2880(1620) ,
  \2346(1256) ,
  \1367(799) ,
  \3112(1464) ,
  \2512(1314) ,
  \1755(225) ,
  \1258(674) ,
  \3069(1073) ,
  \3082(165) ,
  \1069(311) ,
  \2874(129) ,
  \2079(745) ,
  \1924(791) ,
  \2827(1630) ,
  \678(275) ,
  \1006(409) ,
  \3379(1478) ,
  \3369(1477) ,
  \1409(917) ,
  \2966(220) ,
  \1030(1442) ,
  \2854(1685) ,
  \1307(954) ,
  \1418(769) ,
  \1433(636) ,
  \917(549) ,
  \1060(243) ,
  \717(120) ,
  \1603(1031) ,
  \1356(906) ,
  \2519(1300) ,
  \1487(844) ,
  \1666(1133) ,
  \3272(1262) ,
  \938(722) ,
  \1323(815) ,
  \3071(1014) ,
  \2202(994) ,
  \3498(1636) ,
  \3366(1364) ,
  \954(1532) ,
  \1600(1087) ,
  \3035(394) ,
  \2681(1574) ,
  \2647(1372) ,
  \3147(1242) ,
  \1342(663) ,
  \1662(1418) ,
  \1437(860) ,
  \1498(624) ,
  \1415(715) ,
  \3170(1045) ,
  \2734(558) ,
  \2371(1199) ,
  \2236(748) ,
  \3465(1505) ,
  \1883(1011) ,
  \460(89) ,
  \1930(936) ,
  \1909(545) ,
  \2603(1488) ,
  \1255(833) ,
  \1243(609) ,
  \617(536) ,
  \2536(1440) ,
  \1756(360) ,
  \788(109) ,
  \3459(1485) ,
  \3013(174) ,
  \1271(827) ,
  \2716(464) ,
  \1453(861) ,
  \1623(1387) ,
  \2931(60) ,
  \897(168) ,
  \1204(517) ,
  \911(724) ,
  \2098(989) ,
  \2062(395) ,
  \907(67) ,
  \1530(302) ,
  \2844(1662) ,
  \2668(1576) ,
  \2272(1182) ,
  \432(99) ,
  \2298(237) ,
  \2495(1283) ,
  \3110(251) ,
  \501(79) ,
  \3513(1613) ,
  \1156(373) ,
  \1834(215) ,
  \932(1371) ,
  \1022(206) ,
  \1618(578) ,
  \2970(491) ,
  \3182(982) ,
  \3166(980) ,
  \981(314) ,
  \2877(217) ,
  \2415(1287) ,
  \2255(987) ,
  \2593(1489) ,
  \2623(1470) ,
  \2210(1107) ,
  \1439(841) ,
  \586(356) ,
  \1405(858) ,
  \1629(566) ,
  \3219(1267) ,
  \1262(706) ,
  \1326(678) ,
  \1353(875) ,
  \802(100) ,
  \569(796) ,
  \3047(546) ,
  \3305(1380) ,
  \1497(608) ,
  \2341(945) ,
  \408(1660) ,
  \649(723) ,
  \1455(842) ,
  \2375(1097) ,
  \1421(859) ,
  \1764(488) ,
  \1072(374) ,
  \1249(806) ,
  \2963(133) ,
  \3531(1691) ,
  \1250(813) ,
  \668(425) ,
  \2358(1196) ,
  \2658(1575) ,
  \492(80) ,
  \901(542) ,
  \1745(187) ,
  \3103(71) ,
  \386(1602) ,
  \2699(569) ,
  \2585(1411) ,
  \1471(843) ,
  \1501(640) ,
  \1534(431) ,
  \2362(1234) ,
  \1282(829) ,
  \903(264) ,
  \1231(511) ,
  \1829(214) ,
  \1856(417) ,
  \2983(359) ,
  \2805(1446) ,
  \2780(1580) ,
  \2670(1551) ,
  \2760(1391) ,
  \1057(197) ,
  \2667(1569) ,
  \2757(1579) ,
  \2150(1102) ,
  \1322(809) ,
  \2021(283) ,
  \1488(778) ,
  \799(101) ,
  \3451(1487) ,
  \3361(1476) ,
  \1407(839) ,
  \1298(644) ,
  \2167(384) ,
  \1397(698) ,
  \1410(667) ,
  \2718(570) ,
  \1277(611) ,
  \1826(123) ,
  \1108(371) ,
  \2004(737) ,
  \759(198) ,
  \2553(1531) ,
  \3302(1348) ,
  \589(880) ,
  \2896(1648) ,
  \1582(1020) ,
  \3497(1554) ,
  \2349(1232) ,
  \2859(1708) ,
  \898(84) ,
  \2313(1209) ,
  \1656(552) ,
  \3130(1201) ,
  \3378(1299) ,
  \3002(971) ,
  \2739(1501) ,
  \3520(1661) ,
  \855(330) ,
  \1676(1282) ,
  \1508(755) ,
  \1542(348) ,
  \3134(986) ,
  \1734(232) ,
  \1605(310) ,
  \1010(326) ,
  \2833(1681) ,
  \2445(1098) ,
  \906(156) ,
  \1423(840) ,
  \1382(633) ,
  \591(965) ,
  \3053(731) ,
  \2511(1313) ,
  \2455(1095) ,
  \2697(463) ,
  \2531(1312) ,
  \2131(746) ,
  \1622(1351) ,
  \2483(999) ,
  \1288(822) ,
  \2660(1584) ,
  \2592(1508) ,
  \2797(1582) ,
  \2007(401) ,
  \2956(224) ,
  \3528(1697) ,
  \2040(996) ,
  \1359(664) ,
  \2526(1370) ,
  \595(837) ,
  \603(1120) ,
  \1735(365) ,
  \1001(203) ,
  \1345(615) ,
  \608(1185) ,
  \707(127) ,
  \3568(1694) ,
  \3102(249) ,
  \2177(846) ,
  \2288(240) ,
  \1029(588) ,
  \2190(922) ,
  \980(200) ,
  \2219(380) ,
  \1496(688) ,
  \1974(743) ,
  \1599(1029) ,
  \3211(1266) ,
  \2579(1450) ,
  \2612(1272) ,
  \3386(1423) ,
  \1889(998) ,
  \1744(298) ,
  \1895(1115) ,
  \1472(779) ,
  \2156(1145) ,
  \1675(1134) ,
  \1602(1030) ,
  \2099(963) ,
  \2937(146) ,
  \1772(212) ,
  \2615(1447) ,
  \701(523) ,
  \483(81) ,
  \1645(581) ,
  \1456(780) ,
  \1016(319) ,
  \3040(152) ,
  \645(890) ,
  \2925(1629) ,
  \2950(55) ,
  \2293(238) ,
  \1732(287) ,
  \3422(1311) ,
  \1615(1263) ,
  \1366(648) ,
  \663(1124) ,
  \3058(522) ,
  \3236(1041) ,
  \1679(1188) ,
  \3245(1172) ,
  \2572(1510) ,
  \550(136) ,
  \545(147) ,
  \2205(1055) ,
  \1740(385) ,
  \2728(1599) ,
  \401(1716) ,
  \986(958) ,
  \1438(851) ,
  \1256(957) ,
  \1871(499) ,
  \1364(712) ,
  \3046(387) ,
  \1291(660) ,
  \3043(254) ,
  \1299(825) ,
  \2672(1524) ,
  \1019(382) ,
  \2544(1400) ,
  \1279(707) ,
  \2939(58) ,
  \1435(763) ,
  \3304(1373) ,
  \1760(291) ,
  \2351(1152) ,
  \3155(1180) ,
  \3517(1672) ,
  \1454(852) ,
  \848(73) ,
  \1400(650) ,
  \1942(1154) ,
  \2320(948) ,
  \1275(675) ,
  \3142(1143) ,
  \1724(184) ,
  \3111(1482) ,
  \1408(783) ,
  \597(960) ,
  \3186(1047) ,
  \1817(459) ,
  \1339(801) ,
  \1470(853) ,
  \2085(928) ,
  \2350(1195) ,
  \904(412) ,
  \1032(115) ,
  \588(137) ,
  \1301(893) ,
  \3185(1217) ,
  \1554(471) ,
  \1659(1386) ,
  \1758(300) ,
  \1450(637) ,
  \571(942) ,
  \3401(1454) ,
  \1426(916) ,
  \982(322) ,
  \3086(263) ,
  \3224(975) ,
  \2953(138) ,
  \1997(1075) ,
  \357(1136) ,
  \2302(236) ,
  \1424(782) ,
  \1324(953) ,
  \3552(1610) ,
  \1933(1117) ,
  \1614(1325) ,
  \2973(591) ,
  \2625(1360) ,
  \1020(398) ,
  \3338(1452) ,
  \2256(959) ,
  \1736(500) ,
  \942(441) ,
  \2400(1192) ,
  \2338(1153) ,
  \1413(619) ,
  \2426(1307) ,
  \928(576) ,
  \2399(1229) ,
  \991(404) ,
  \1427(668) ,
  \352(260) ,
  \2826(1617) ,
  \1527(284) ,
  \807(181) ,
  \2229(836) ,
  \1853(735) ,
  \993(544) ,
  \3138(1051) ,
  \3470(1601) ,
  \2843(1651) ,
  \1440(781) ,
  \2137(925) ,
  \3128(1050) ,
  \3285(1413) ,
  \1672(584) ,
  \3286(1407) ,
  \2662(1548) ,
  \3560(1693) ,
  \2626(1395) ,
  \1284(902) ,
  \2401(1350) ,
  \2424(1277) ,
  \3256(1409) ,
  \1195(507) ,
  \1768(351) ,
  \673(1082) ,
  \1596(1086) ,
  \3079(91) ,
  \2719(1538) ,
  \823(180) ,
  \2387(1190) ,
  \442(98) ,
  \2733(465) ,
  \1535(422) ,
  \2853(1652) ,
  \3240(977) ,
  \3502(1628) ,
  \3433(1529) ,
  \3235(1211) ,
  \1422(850) ,
  \3124(985) ,
  \3154(1168) ,
  \1399(634) ,
  \685(427) ,
  \1412(603) ,
  \1922(478) ,
  \1272(830) ,
  \2474(930) ,
  \2539(1480) ,
  \2022(489) ,
  \2242(919) ,
  \831(92) ,
  \2599(1527) ,
  \1300(883) ,
  \2372(1203) ,
  \2607(1301) ,
  \1591(1025) ,
  \1159(510) ,
  \1386(888) ,
  \1370(866) ,
  \2552(1546) ,
  \2666(1565) ,
  \2031(932) ,
  \1432(716) ,
  \956(346) ,
  \1489(771) ,
  \3398(1332) ,
  \1671(1358) ,
  \607(1158) ,
  \2725(1389) ,
  \700(1160) ,
  \1355(896) ,
  \1670(1225) ,
  \2803(562) ,
  \1343(679) ,
  \553(227) ,
  \1021(529) ,
  \2478(64) ,
  \2999(974) ,
  \1048(62) ,
  \1075(512) ,
  \1619(447) ,
  \2634(1416) ,
  \3264(1384) ,
  \3284(1382) ,
  \1624(1318) ,
  \2964(131) ,
  \2114(388) ,
  \1147(508) ,
  \3516(1650) ,
  \1585(305) ,
  \3458(1455) ,
  \2788(1503) ,
  \1726(396) ,
  \3077(1074) ,
  \2584(1437) ,
  \1723(295) ,
  \1870(280) ,
  \839(78) ,
  \3308(1260) ,
  \3006(1037) ,
  \1312(693) ,
  \3395(1429) ,
  \3482(1665) ,
  \951(1564) ,
  \3387(1479) ,
  \1431(700) ,
  \2517(1302) ,
  \3557(1695) ,
  \3298(1316) ,
  \2500(1319) ,
  \2146(1108) ,
  \983(908) ,
  \1294(612) ,
  \1791(344) ,
  \1827(122) ,
  \1251(819) ,
  \3195(1235) ,
  \2832(1674) ,
  \1541(151) ,
  \2431(1226) ,
  \2525(1377) ,
  \1598(1028) ,
  \2010(537) ,
  \3418(1331) ,
  \2309(1206) ,
  \1646(436) ,
  \696(429) ,
  \2523(1200) ,
  \2608(1339) ,
  \2216(740) ,
  \3116(1494) ,
  \610(432) ,
  \583(1094) ,
  \702(530) ,
  \1750(494) ,
  \2735(571) ,
  \392(1594) ,
  \1509(752) ,
  \1084(375) ,
  \400(1715) ,
  \2892(1678) ,
  \2564(1435) ,
  \1643(727) ,
  \2041(990) ,
  \3354(1365) ,
  \1790(194) ,
  \1616(733) ,
  \2164(739) ,
  \1035(63) ,
  \1417(651) ,
  \1457(773) ,
  \3267(1460) ,
  \2091(1008) ,
  \1812(458) ,
  \530(66) ,
  \1996(1062) ,
  \1354(886) ,
  \3549(1633) ,
  \3443(1507) ,
  \2518(1274) ,
  \929(734) ,
  \3205(1239) ,
  \1473(772) ,
  \1763(358) ,
  \988(315) ,
  \3030(161) ,
  \990(267) ,
  \1467(638) ,
  \1049(114) ,
  \2157(1169) ,
  \2059(738) ,
  \2571(1473) ,
  \2581(1472) ,
  \1411(683) ,
  \2601(1471) ,
  \3033(258) ,
  \916(442) ,
  \1320(904) ,
  \2181(277) ,
  \570(798) ,
  \1874(792) ,
  \1500(720) ,
  \1762(223) ,
  \1013(403) ,
  \944(969) ,
  \1317(873) ,
  \2370(1236) ,
  \1350(807) ,
  \1376(665) ,
  \2268(1245) ,
  \3109(159) ,
  \2849(1673) ,
  \1859(547) ,
  \1289(826) ,
  \2530(1141) ,
  \3489(1656) ,
  \2960(52) ,
  \2475(927) ,
  \2920(1711) ,
  \2638(1483) ,
  \1673(439) ,
  \3095(72) ,
  \2076(279) ,
  \1043(149) ,
  \1916(1077) ,
  \689(1125) ,
  \1425(775) ,
  \2124(1070) ,
  \672(533) ,
  \2633(1420) ,
  \2938(144) ,
  \1880(938) ,
  \864(210) ,
  \867(332) ,
  \389(1592) ,
  \902(729) ,
  \1246(625) ,
  \1429(604) ,
  \3350(1334) ,
  \3454(1432) ,
  \395(1486) ,
  \2578(1511) ,
  \721(211) ,
  \1362(616) ,
  \2170(525) ,
  \2111(1035) ,
  \3499(1540) ,
  \3119(1518) ,
  \1383(649) ,
  \1441(774) ,
  \640(541) ,
  \724(119) ,
  \2025(789) ,
  \1443(915) ,
  \3253(1352) ,
  \1452(758) ,
  \2233(278) ,
  \680(420) ,
  \1449(717) ,
  \1609(577) ,
  \2317(1156) ,
  \1273(956) ,
  \1381(713) ,
  \2913(1688) ,
  \642(262) ,
  \2017(872) ,
  \2289(239) ,
  \3410(1330) ,
  \356(1135) ,
  \1972(493) ,
  \1268(812) ,
  \1005(392) ,
  \2994(970) ,
  \3301(1306) ,
  \1017(327) ,
  \1242(593) ,
  \1296(708) ,
  \1038(148) ,
  \2538(1481) ,
  \551(134) ,
  \3276(1292) ,
  \2541(1498) ,
  \826(96) ,
  \546(145) ,
  \1954(736) ,
  \1590(1024) ,
  \565(795) ,
  \3290(1315) ,
  \3446(1495) ,
  \1014(962) ,
  \943(445) ,
  \1384(784) ,
  \3362(1398) ,
  \3382(1396) ,
  \3208(1139) ,
  \1361(600) ,
  \1329(694) ,
  \3466(1606) ,
  \1000(538) ,
  \2675(1562) ,
  \2490(1230) ,
  \2203(988) ,
  \2391(944) ,
  \362(1441) ,
  \1374(907) ,
  \1008(204) ,
  \2128(276) ,
  \2555(1566) ,
  \3280(1349) ,
  \1680(1359) ,
  \860(208) ,
  \1448(701) ,
  \3541(1632) ,
  \2954(135) ,
  \2484(1052) ,
  \1341(952) ,
  \3449(1525) ,
  \2043(1059) ,
  \2665(1558) ,
  \2540(1462) ,
  \845(74) ,
  \3330(1310) ,
  \2567(1333) ,
  \1292(676) ,
  \2524(1375) ,
  \1537(1018) ,
  \616(424) ,
  \1752(188) ,
  \2357(1233) ,
  \987(201) ,
  \1387(877) ,
  \1444(669) ,
  \2752(559) ,
  \2222(520) ,
  \3442(1519) ,
  \1026(354) ,
  \3005(1039) ,
  \1886(1005) ,
  \567(941) ,
  \3283(1376) ,
  \3536(1698) ,
  \1739(288) ,
  \3475(1641) ,
  \1120(376) ,
  \2173(845) ,
  \2679(555) ,
  \3548(1621) ,
  \2548(1530) ,
  \2433(1251) ,
  \2182(483) ,
  \1990(997) ,
  \2694(1612) ,
  \3394(1424) ,
  \1828(110) ,
  \3293(1379) ,
  \3066(1066) ,
  \2771(1523) ,
  \1747(381) ,
  \1018(253) ,
  \1719(402) ,
  \576(793) ,
  \2278(207) ,
  \1647(551) ,
  \1267(805) ,
  \1430(620) ,
  \1261(690) ,
  \3441(1543) ,
  \3334(1426) ,
  \2485(369) ,
  \998(397) ,
  \3339(1517) ,
  \1314(629) ,
  \3054(726) ,
  \2558(1493) ,
  \1771(485) ,
  \2967(497) ,
  \2598(1490) ,
  \1538(548) ,
  \2557(1451) ,
  \582(1092) ,
  \2921(1701) ,
  \1890(992) ,
  \1428(684) ,
  \1511(911) ,
  \3406(1297) ,
  \3244(1042) ,
  \2802(469) ,
  \1587(1023) ,
  \1927(935) ,
  \2103(1110) ,
  \2617(1469) ,
  \1741(230) ,
  \2838(1682) ,
  \2748(1522) ,
  \1504(777) ,
  \1894(1078) ,
  \758(108) ,
  \3481(1655) ,
  \870(443) ,
  \2052(213) ,
  \3204(1049) ,
  \3287(1346) ,
  \2537(1463) ,
  \1767(292) ,
  \3085(172) ,
  \456(94) ,
  \1971(282) ,
  \2831(1664) ,
  \1025(244) ,
  \3163(1181) ,
  \1469(754) ,
  \360(794) ,
  \2597(1509) ,
  \1310(597) ,
  \2199(1001) ,
  \989(323) ,
  \1027(393) ,
  \1901(336) ,
  \2023(476) ,
  \1340(808) ,
  \1371(876) ,
  \2077(487) ,
  \3020(163) ,
  \2234(480) ,
  \1742(364) ,
  \1360(680) ,
  \1617(1356) ,
  \1283(892) ,
  \1597(308) ,
  \1902(451) ,
  \2891(1669) ,
  \2143(1116) ,
  \3277(1345) ,
  \3491(1539) ,
  \804(303) ,
  \540(65) ,
  \1490(765) ,
  \2871(128) ,
  \794(182) ,
  \1612(1127) ,
  \1458(767) ,
  \1252(824) ,
  \1244(689) ,
  \3194(1048) ,
  \554(219) ,
  \3007(97) ,
  \3326(1279) ,
  \[10] ,
  \1636(580) ,
  \2978(492) ,
  \2622(1422) ,
  \3212(1163) ,
  \1379(617) ,
  \[11] ,
  \1066(312) ,
  \2037(1003) ,
  \2225(835) ,
  \1087(514) ,
  \1304(810) ,
  \1398(714) ,
  \[12] ,
  \1604(1088) ,
  \1620(565) ,
  \1751(299) ,
  \[13] ,
  \643(413) ,
  \1334(864) ,
  \3346(1453) ,
  \3419(51) ,
  \3078(1121) ,
  \[14] ,
  \3193(1212) ,
  \3150(1144) ,
  \2129(484) ,
  \2204(961) ,
  \933(1419) ,
  \1607(1033) ,
  \1474(766) ,
  \1941(1123) ,
  \1674(554) ,
  \714(124) ,
  \2345(1194) ,
  \681(1081) ,
  \1319(894) ,
  \1434(652) ,
  \3023(268) ,
  \[17] ,
  \2065(534) ,
  \3034(255) ,
  \[18] ,
  \3385(1496) ,
  \2476(924) ,
  \[19] ,
  \661(1080) ,
  \619(1091) ,
  \3563(1702) ,
  \2577(1474) ,
  \3025(406) ,
  \1028(521) ,
  \2562(1410) ,
  \3510(1625) ,
  \1633(1257) ,
  \3478(1653) ,
  \2409(1285) ,
  \2354(946) ,
  \1368(847) ,
  \1957(407) ,
  \1259(594) ,
  \1987(1004) ,
  \3434(1552) ,
  \2439(1281) ,
  \1975(790) ,
  \2888(1668) ,
  \3010(173) ,
  \2769(560) ,
  \2251(1000) ,
  \1632(1326) ,
  \2848(1663) ,
  \665(433) ,
  \1626(1417) ,
  \1378(601) ,
  \1484(639) ,
  \2600(1542) ,
  \1023(320) ,
  \3402(1361) ,
  \2570(1491) ,
  \978(379) ,
  \[20] ,
  \2632(1415) ,
  \851(68) ,
  \1096(370) ,
  \[21] ,
  \836(85) ,
  \3331(1516) ,
  \3203(1213) ,
  \1545(470) ,
  \1998(1112) ,
  \2331(1294) ,
  \2916(1712) ,
  \1799(461) ,
  \3525(1686) ,
  \397(1394) ,
  \349(1224) ,
  \2395(1191) ,
  \3426(1344) ,
  \2736(1502) ,
  \2419(1288) ,
  \2645(1305) ,
  \1358(951) ,
  \3036(400) ,
  \1731(185) ,
  \3090(166) ,
  \1186(505) ,
  \1584(1083) ,
  \3565(1696) ,
  \2774(1572) ,
  \1303(803) ,
  \2700(1520) ,
  \2942(57) ,
  \1392(918) ,
  \447(95) ,
  \2804(575) ,
  \1718(285) ,
  \398(1366) ,
  \1765(301) ,
  \635(164) ,
  \2677(1514) ,
  \1442(768) ,
  \566(797) ,
  \2117(531) ,
  \1721(368) ,
  \1502(656) ,
  \3055(532) ,
  \1663(583) ,
  \3490(1667) ,
  \2974(589) ,
  \2909(1684) ,
  \1318(884) ,
  \1290(955) ,
  \941(333) ,
  \1447(621) ,
  \1757(490) ,
  \596(854) ,
  \1278(691) ,
  \2563(1378) ,
  \2332(1264) ,
  \3158(979) ,
  \1536(1016) ,
  \1720(235) ,
  \2794(1392) ,
  \1510(750) ,
  \2586(1459) ,
  \1446(605) ,
  \3213(1240) ,
  \1981(934) ,
  \2823(1631) ,
  \2554(1560) ,
  \1872(479) ,
  \1393(666) ,
  \1388(867) ,
  \1581(304) ,
  \657(177) ,
  \552(132) ,
  \547(143) ,
  \1063(242) ,
  \2185(786) ,
  \741(116) ,
  \1054(196) ,
  \1862(899) ,
  \3120(1513) ,
  \2602(1449) ,
  \1460(914) ,
  \1466(718) ,
  \3037(157) ,
  \3316(1341) ,
  \3026(410) ,
  \2359(1258) ,
  \887(444) ,
  \2754(1556) ,
  \2072(863) ,
  \2248(1006) ,
  \479(82) ,
  \979(543) ,
  \1357(800) ,
  \2333(1317) ,
  \605(1186) ,
  \3190(983) ,
  \3174(981) ,
  \1263(626) ,
  \1327(598) ,
  \1769(221) ,
  \3275(1461) ,
  \861(209) ,
  \2533(1193) ,
  \2155(1150) ,
  \2379(1250) ,
  \1050(113) ,
  \2547(1545) ,
  \2237(785) ,
  \2765(1590) ,
  \1586(1022) ,
  \1730(296) ,
  \2868(50) ,
  \2860(1710) ,
  \1346(695) ,
  \3403(1402) ,
  \1947(1170) ,
  \950(1547) ,
  \1661(1126) ,
  \2751(466) ,
  \1269(818) ,
  \2042(964) ,
  \3259(1383) ,
  \736(118) ,
  \1465(702) ,
  \1377(681) ,
  \2678(462) ,
  \560(226) ,
  \1002(317) ,
  \590(891) ,
  \3070(1119) ,
  \1939(1105) ,
  \3179(1179) ,
  \1123(516) ,
  \1639(1130) ,
  \1111(506) ,
  \1613(1293) ,
  \654(256) ,
  \3494(1627) ,
  \3337(1534) ,
  \704(126) ,
  \3547(1645) ,
  \997(259) ,
  \3524(1671) ,
  \3438(1500) ,
  \2102(1071) ,
  \555(231) ,
  \2837(1675) ,
  \1247(641) ,
  \2917(1703) ,
  \780(106) ,
  \2285(241) ,
  \2209(1068) ,
  \1007(528) ,
  \3532(1705) ,
  \1621(1128) ,
  \2680(568) ,
  \992(418) ,
  \1177(515) ,
  \2386(1227) ,
  \1461(670) ,
  \1991(991) ,
  \3319(1367) ,
  \1960(540) ,
  \562(363) ,
  \1681(192) ,
  \1601(309) ,
  \3355(1457) ,
  \2505(1320) ,
  \1794(460) ,
  \1893(1064) ,
  \3430(1537) ,
  \557(366) ,
  \3216(1140) ,
  \1338(905) ,
  \1402(889) ,
  \3329(1162) ,
  \3572(1700) ,
  \641(728) ,
  \1445(685) ,
  \1606(1032) ,
  \3474(1618) ,
  \2183(473) ,
  \3229(1174) ,
  \842(77) ,
  \2378(1278) ,
  \2308(1271) ,
  \2028(931) ,
  \354(257) ,
  \995(316) ,
  \1642(1259) ,
  \1459(762) ,
  \1373(897) ,
  \2663(1567) ,
  \1331(630) ,
  \2986(355) ,
  \1132(377) ,
  \625(167) ,
  \1637(449) ,
  \913(390) ,
  \2816(1468) ,
  \2556(1475) ,
  \1505(770) ,
  \1641(1327) ,
  \2013(871) ,
  \3050(539) ,
  \3145(1268) ,
  \1475(761) ,
  \1748(228) ,
  \634(247) ,
  \1351(855) ,
  \1722(502) ,
  \1222(509) ,
  \1315(645) ,
  \579(939) ,
  \1770(357) ,
  \2703(1578) ,
  \1308(661) ,
  \1923(742) ,
  \1414(699) ,
  \2908(1676) ,
  \3024(261) ,
  \3370(1399) ,
  \1390(848) ,
  \1610(446) ,
  \1486(751) ,
  \2080(788) ,
  \3409(1430) ,
  \2900(350) ,
  \1011(909) ,
  \1240(657) ,
  \1759(189) ,
  \1491(760) ,
  \2003(453) ,
  \976(266) ,
  \3390(1397) ,
  \1754(353) ,
  \2929(1644) ,
  \1664(438) ,
  \3564(1699) ,
  \671(426) ,
  \604(1159) ,
  \2078(475) ,
  \1396(618) ,
  \2684(1596) ,
  \3462(1593) ,
  \2235(472) ,
  \1634(730) ,
  \2763(1589) ,
  \2998(1036) ,
  \2609(1369) ,
  \2821(1607) ,
  \2673(1557) ,
  \2945(142) ,
  \2808(1443) ,
  \2535(1338) ,
  \731(121) ,
  \2989(486) ,
  \915(331) ,
  \1984(1010) ,
  \2753(572) ,
  \2152(1149) ,
  \662(550) ,
  \1477(913) ,
  \636(175) ,
  \1253(828) ,
  \3248(978) ,
  \2425(1249) ,
  \791(103) ,
  \3171(1178) ,
  \1372(887) ,
  \2852(1639) ,
  \1669(1252) ,
  \1451(653) ,
  \1305(816) ,
  \2477(921) ,
  \2002(338) ,
  \2635(1465) ,
  \655(416) ,
  \3450(1515) ,
  \1668(1323) ,
  \2315(1244) ,
  \890(125) ,
  \526(69) ,
  \2193(923) ,
  \363(1466) ,
  \1031(1571) ,
  \3295(1276) ,
  \1660(1308) ,
  \1276(595) ,
  \1395(602) ,
  \3243(1207) ,
  \3014(271) ,
  \1595(1027) ,
  \2713(1588) ,
  \2458(1096) ,
  \1967(882) ,
  \3074(1067) ,
  \3483(1642) ,
  \1335(874) ,
  \2101(1058) ,
  \2786(561) ,
  \1389(857) ,
  \2254(993) ,
  \3342(1427) ,
  \2842(1638) ,
  \2097(995) ,
  \2491(1255) ,
  \2768(467) ,
  \3556(1622) ,
  \2132(787) ,
  \1024(328) ,
  \2576(1492) ,
  \2981(592) ,
  \3427(1512) ,
  \2261(1065) ,
  \620(1093) ,
  \644(269) ,
  \1572(334) ,
  \2621(1448) ,
  \1419(879) ,
  \3169(1220) ,
  \3094(265) ,
  \2265(1215) ,
  \3131(1184) ,
  \3121(1183) ,
  \3221(1173) ,
  \1375(950) ,
  \3016(419) ,
  \2650(1404) ,
  \660(274) ,
  \1248(834) ,
  \1635(1355) ,
  \2589(1362) ,
  \994(202) ,
  \3414(1298) ,
  \2275(1246) ,
  \1015(205) ,
  \2448(1099) ,
  \2514(1309) ,
  \1540(111) ,
  \3027(162) ,
  \1295(692) ,
  \3269(1439) ,
  \3320(1374) ,
  \2629(1385) ,
  \690(535) ,
  \1749(362) ,
  \3113(1499) ,
  \1993(1061) ,
  \2928(1623) ,
  \639(272) ,
  \1464(622) ,
  \3252(1043) ,
  \3506(1637) ,
  \1478(671) ,
  \2482(949) ,
  \548(141) ,
  \614(968) ,
  \1651(1261) ,
  \2088(929) ,
  \974(313) ,
  \1648(1131) ,
  \2451(1142) ,
  \3457(1506) ,
  \3232(976) ,
  \1213(519) ,
  \1316(820) ,
  \2245(920) ,
  \1973(477) ,
  \2676(1533) ,
  \1746(289) ,
  \1877(937) ,
  \3061(725) ,
  \2461(1137) ,
  \1630(1129) ,
  \3129(1237) ,
  \1627(579) ,
  \833(86) ,
  \669(1019) ,
  \3161(1219) ,
  \3322(1401) ,
  \1483(719) ,
  \1512(193) ,
  \513(75) ,
  \1593(307) ,
  \2624(1329) ,
  \1658(1342) ,
  \1638(567) ,
  \1891(967) ,
  \3358(1363) ,
  \3374(1273) ,
  \1348(631) ,
  \3063(1013) ,
  \3507(1598) ,
  \1738(186) ,
  \568(972) ,
  \893(216) ,
  \1892(1063) ,
  \2501(1353) ,
  \1051(112) ,
  \3220(1164) ,
  \404(1714) ,
  \1286(811) ,
  \1280(627) ,
  \2363(1197) ,
  \3139(1241) ,
  \2865(61) ,
  \2481(150) ,
  \1344(599) ,
  \2822(1619) ,
  \3162(1044) ,
  \2151(1122) ,
  \2271(1114) ,
  \2307(1270) ,
  \350(1223) ,
  \1463(606) ,
  \679(1015) ,
  \2922(1608) ,
  \3571(1704) ,
  \3486(1654) ,
  \2489(1100) ,
  \2262(1106) ,
  \1394(682) ,
  \3393(1497) ,
  \3106(154) ,
  \561(229) ,
  \2047(1072) ,
  \2130(474) ,
  \1403(878) ,
  \1650(1322) ,
  \2364(1151) ,
  \1766(190) ,
  \1482(703) ,
  \2068(862) ,
  \973(199) ,
  \1852(450) ,
  \3523(1680) ,
  \1936(1113) ,
  \476(83) ,
  \1945(1155) ,
  \923(482) ,
  \1257(658) ,
  \2208(1056) ,
  \2910(1689) ,
  \606(1118) ,
  \2444(1166) ,
  \2454(1165) ,
  \688(428) ,
  \2839(1614) ,
  \1003(325) ,
  \947(910) ,
  \517(70) ,
  \2534(1335) ,
  \977(414) ,
  \996(324) ,
  \1264(642) ,
  \556(233) ,
  \1592(1085) ,
  \1649(1291) ,
  \2464(1248) ,
  \2864(1709) ,
  \2024(744) ,
  \1416(635) ,
  \3533(1687) ,
  \2344(1231) ,
  \2388(1147) ,
  \1728(367) ,
  \1727(234) ,
  \806(293) ,
  \1468(654) ,
  \1506(764) ,
  \1851(335) ,
  \366(1577) ,
  \1285(804) ,
  \1906(411) ,
  \1665(553) ,
  \3200(984) ,
  \1363(696) ,
  \380(1615) ,
  \2527(1412) ,
  \1611(564) ,
  \1391(838) ,
  \2836(1666) ,
  \1631(1286) ;
assign
  \703(1187)  = \702(530)  | (\701(523)  | \700(1160) ),
  \2580(1425)  = ~\3378(1299)  | ~\3371(1405) ,
  \920(361)  = \915(331)  & \588(137) ,
  \2886(1658)  = ~\3547(1645)  | ~\3544(1609) ,
  \2742(1390)  = \2735(571)  & \1644(1354) ,
  \2997(1038)  = ~\2991(973) ,
  \574(585)  = ~\2989(486)  | ~\2986(355) ,
  \1539(1079)  = \1538(548)  | (\1537(1018)  | \1536(1016) ),
  \2907(1683)  = \2903(349)  & (\2892(1678)  & \2844(1662) ),
  \1476(757)  = \1468(654)  & \317(42) ,
  \699(430)  = \806(293)  & \804(303) ,
  \3261(1438)  = \2527(1412) ,
  \912(250)  = ~\3109(159)  | ~\3106(154) ,
  \1678(1254)  = ~\2400(1192)  | ~\2399(1229) ,
  \3196(1198)  = ~\3194(1048)  | ~\3187(1176) ,
  \2325(1204)  = \1947(1170) ,
  \1940(1103)  = \1927(935)  & (\1916(1077)  & \200(25) ),
  \2782(1581)  = ~\2777(1445)  & (~\2774(1572)  & ~\2771(1523) ),
  \3473(1604)  = ~\3467(1591) ,
  \3268(1414)  = ~\3264(1384) ,
  \2654(1337)  = \2519(1300) ,
  \776(107)  = \33(3) ,
  \1677(1324)  = \1673(439)  & \1676(1282) ,
  \2659(1568)  = \2638(1483)  & (\2549(1559)  & (\2558(1493)  & \2572(1510) )),
  \463(88)  = ~\68(8) ,
  \1135(518)  = \1132(377) ,
  \784(191)  = \780(106) ,
  \2730(1600)  = ~\2725(1389)  & (~\2722(1586)  & ~\2719(1538) ),
  \1733(389)  = \1730(296)  & \97(11) ,
  \2903(349)  = ~\2897(49)  | ~\2877(217) ,
  \2467(1275)  = \2464(1248) ,
  \910(527)  = ~\913(390)  | ~\912(250) ,
  \1492(756)  = \1484(639)  & \317(42) ,
  \1594(1026)  = \1593(307)  & \1324(953) ,
  \387(1616)  = \[12] ,
  \2722(1586)  = \2717(557)  & \2668(1576) ,
  \2991(973)  = \571(942) ,
  \2162(341)  = ~\1834(215) ,
  \1144(372)  = ~\1063(242)  | ~\1038(148) ,
  \1737(297)  = ~\1681(192) ,
  \985(378)  = \982(322)  & \159(21) ,
  \2100(1057)  = \2094(1002)  | \2091(1008) ,
  \1725(286)  = \1699(105)  & \1681(192) ,
  \2947(56)  = \250(33) ,
  \1325(662)  = ~\1075(512) ,
  \1009(318)  = ~\759(198) ,
  \1270(823)  = \1262(706)  & \137(18) ,
  \2336(1295)  = ~\3153(1269)  | ~\3150(1144) ,
  \2828(1640)  = ~\2827(1630)  | ~\2826(1617) ,
  \896(176)  = ~\45(5)  | (~\732(117)  | ~\717(120) ),
  \1311(613)  = ~\1111(506) ,
  \3411(1403)  = \2609(1369) ,
  \648(526)  = ~\647(391)  | ~\646(248) ,
  \2669(1563)  = ~\3441(1543)  | ~\3438(1500) ,
  \2549(1559)  = ~\2548(1530)  | ~\2547(1545) ,
  \2274(1214)  = ~\1895(1115)  | (~\1998(1112)  | (~\1947(1170)  | ~\2043(1059) )),
  \1004(252)  = \1001(203)  & \906(156) ,
  \650(273)  = \621(170)  & \432(99) ,
  \504(76)  = \97(11) ,
  \927(347)  = ~\893(216) ,
  \1462(686)  = ~\1177(515) ,
  \1385(898)  = \1377(681)  & \447(95) ,
  \2196(1007)  = \2190(922)  & (\2173(845)  & \169(22) ),
  \[0]  = ~\352(260) ,
  \2488(503)  = ~\2485(369) ,
  \2965(218)  = ~\2963(133)  | ~\2960(52) ,
  \2717(557)  = ~\870(443) ,
  \2149(1104)  = \2140(926)  & (\2124(1070)  & \190(24) ),
  \[1]  = ~\354(257) ,
  \3515(1635)  = ~\3513(1613)  | ~\3510(1625) ,
  \[2]  = ~\360(794)  | ~\359(587) ,
  \2140(926)  = ~\2132(787) ,
  \1644(1354)  = ~\1643(727)  & (~\1641(1327)  & ~\1639(1130) ),
  \1654(582)  = ~\1554(471) ,
  \1652(1090)  = \1647(551)  & \618(1017) ,
  \2745(1521)  = \2742(1390)  | (\2739(1501)  | \2736(1502) ),
  \[3]  = ~\357(1136)  | ~\356(1135) ,
  \1245(705)  = ~\1135(518) ,
  \2214(342)  = ~\1834(215) ,
  \626(158)  = ~\526(69)  | ~\513(75) ,
  \2777(1445)  = \2770(573)  & \1662(1418) ,
  \[4]  = ~\350(1223)  | ~\349(1224) ,
  \1753(290)  = \1699(105)  & \1681(192) ,
  \2163(456)  = \1773(345)  & \1834(215) ,
  \1352(865)  = \1344(599)  & \492(80) ,
  \[5]  = \2265(1215)  & \2309(1206) ,
  \3017(169)  = \463(88) ,
  \3294(1347)  = ~\3290(1315) ,
  \[6]  = ~\368(1296) ,
  \613(423)  = \806(293)  & \804(303) ,
  \[7]  = \398(1366)  | \397(1394) ,
  \1337(895)  = \1329(694)  & \447(95) ,
  \2337(1265)  = ~\3154(1168)  | ~\3147(1242) ,
  \2946(140)  = ~\2942(57) ,
  \[8]  = \363(1466)  & \362(1441) ,
  \1332(646)  = ~\1159(510) ,
  \383(1541)  = ~\2748(1522) ,
  \[9]  = \395(1486)  & \2814(1467) ,
  \3187(1176)  = \2364(1151) ,
  \1266(901)  = \1258(674)  & \432(99) ,
  \2799(1583)  = ~\2794(1392)  & (~\2791(1573)  & ~\2788(1503) ),
  \955(1536)  = ~\3120(1513)  | ~\3113(1499) ,
  \1903(1034)  = \1901(336)  & \986(958) ,
  \467(87)  = \68(8) ,
  \2770(573)  = \870(443)  & \956(346) ,
  \2709(1587)  = \2706(1444)  | (\2703(1578)  | \2700(1520) ),
  \1494(912)  = ~\1493(753)  & (~\1492(756)  & (~\1491(760)  & (~\1490(765)  & (~\1489(771)  & (~\1488(778)  & (~\1487(844)  & ~\1486(751) )))))),
  \1254(831)  = \1246(625)  & \128(16) ,
  \3197(1177)  = \2364(1151) ,
  \1717(183)  = ~\1699(105) ,
  \3015(270)  = ~\3013(174)  | ~\3010(173) ,
  \646(248)  = ~\3101(160)  | ~\3098(153) ,
  \2058(454)  = \1773(345)  & \1834(215) ,
  \1866(900)  = ~\1859(547)  & (~\1856(417)  & ~\1853(735) ),
  \1306(821)  = \1298(644)  & \137(18) ,
  \1330(710)  = ~\1135(518) ,
  \732(117)  = ~\20(2) ,
  \3425(130)  = ~\3419(51) ,
  \2120(1069)  = \2117(531)  | (\2114(388)  | \2111(1035) ),
  \1533(421)  = ~\1527(284) ,
  \2934(59)  = \232(30) ,
  \999(415)  = \996(324)  & \828(93) ,
  \2260(1054)  = ~\2251(1000)  & ~\2248(1006) ,
  \1241(673)  = ~\1087(514) ,
  \3345(1535)  = ~\3339(1517) ,
  \3555(1646)  = ~\3549(1633) ,
  \1921(495)  = \1920(281)  & (\232(30)  & \1817(459) ),
  \2380(1148)  = \2210(1107) ,
  \368(1296)  = \2308(1271)  & \2307(1270) ,
  \984(408)  = \981(314)  & \833(86) ,
  \1297(628)  = ~\1147(508) ,
  \683(434)  = ~\804(303) ,
  \1699(105)  = \33(3)  | \1698(48) ,
  \1309(677)  = ~\1087(514) ,
  \2855(1679)  = ~\3524(1671)  | ~\3517(1672) ,
  \2883(1595)  = \2871(128)  & \2709(1587) ,
  \2643(1328)  = \2642(1304)  & (\2491(1255)  & \330(46) ),
  \1436(870)  = \1428(684)  & \492(80) ,
  \1657(1132)  = \1654(582)  & \1600(1087) ,
  \3505(1555)  = ~\3499(1540) ,
  \2785(468)  = ~\956(346) ,
  \1333(814)  = \1325(662)  & \143(19) ,
  \2508(1381)  = \2419(1288)  & (\2409(1285)  & (\2401(1350)  & \2495(1283) )),
  \3087(90)  = \58(7) ,
  \390(1603)  = \[14] ,
  \1499(704)  = ~\1204(517) ,
  \1912(1076)  = \1909(545)  | (\1906(411)  | \1903(1034) ),
  \3353(1456)  = ~\3347(1434) ,
  \1729(501)  = \1728(367)  | (\1727(234)  | \1726(396) ),
  \2383(943)  = \2173(845)  & \2298(237) ,
  \975(321)  = \759(198)  & \741(116) ,
  \403(1713)  = ~\2921(1701)  | ~\2920(1711) ,
  \828(93)  = \58(7) ,
  \2394(1228)  = ~\3243(1207)  | ~\3240(977) ,
  \1321(802)  = \1313(709)  & \159(21) ,
  \2057(339)  = ~\1834(215) ,
  \2215(457)  = \1773(345)  & \1834(215) ,
  \2982(590)  = ~\2978(492) ,
  \3363(1458)  = \2564(1435) ,
  \3347(1434)  = ~\3286(1407)  | ~\3285(1413) ,
  \3153(1269)  = ~\3147(1242) ,
  \2109(340)  = ~\1834(215) ,
  \3321(1406)  = ~\3319(1367)  | ~\3316(1341) ,
  \3371(1405)  = ~\3304(1373)  | ~\3303(1340) ,
  \1946(1146)  = \1941(1123)  | (\1940(1103)  | \1939(1105) ),
  \3311(1408)  = ~\3305(1380) ,
  \2094(1002)  = \2088(929)  & (\2068(862)  & \179(23) ),
  \926(563)  = ~\887(444) ,
  \2311(1109)  = ~\2100(1057) ,
  \3228(1040)  = ~\3224(975) ,
  \1265(832)  = \1257(658)  & \125(15) ,
  \618(1017)  = \617(536)  | (\616(424)  | \614(968) ),
  \2367(947)  = \2068(862)  & \2289(239) ,
  \1293(596)  = ~\1099(504) ,
  \3237(1171)  = \2388(1147) ,
  \406(1643)  = \2925(1629)  & \2922(1608) ,
  \2930(1649)  = ~\2929(1644)  & ~\2928(1623) ,
  \409(1670)  = \[19] ,
  \2814(1467)  = \2811(1393)  | (\2808(1443)  | \2805(1446) ),
  \3544(1609)  = \2883(1595) ,
  \2034(1009)  = \2028(931)  & (\2013(871)  & \169(22) ),
  \1336(885)  = \1328(614)  & \467(87) ,
  \3540(1706)  = ~\3536(1698) ,
  \2406(1284)  = \2346(1256) ,
  \621(170)  = ~\463(88)  | ~\456(94) ,
  \3062(721)  = ~\3058(522) ,
  \3098(153)  = \907(67) ,
  \1503(749)  = \1495(672)  & \329(45) ,
  \3101(160)  = ~\3095(72) ,
  \1773(345)  = \1772(212)  | \1(0) ,
  \1481(623)  = ~\1195(507) ,
  \1495(672)  = ~\1168(513) ,
  \1404(868)  = \1396(618)  & \492(80) ,
  \1507(759)  = \1499(704)  & \311(41) ,
  \816(179)  = \791(103)  & (\799(101)  & \714(124) ),
  \2257(1053)  = \2251(1000)  | \2248(1006) ,
  \694(435)  = ~\804(303) ,
  \2906(1677)  = \2900(350)  & (\2888(1668)  & \2844(1662) ),
  \2791(1573)  = \2786(561)  & \2675(1562) ,
  \3178(1046)  = ~\3174(981) ,
  \3377(1433)  = ~\3371(1405) ,
  \2863(1707)  = ~\3531(1691)  | ~\3528(1697) ,
  \1168(513)  = \1072(374) ,
  \2594(1526)  = ~\2593(1489)  | ~\2592(1508) ,
  \2661(1561)  = ~\2650(1404)  & ~\2600(1542) ,
  \549(139)  = ~\492(80)  | ~\250(33) ,
  \1313(709)  = ~\1135(518) ,
  \798(102)  = \45(5)  | \41(4) ,
  \1420(869)  = \1412(603)  & \492(80) ,
  \1099(504)  = \1096(370) ,
  \2657(1368)  = ~\2654(1337) ,
  \3177(1216)  = ~\3171(1178) ,
  \692(1157)  = \691(524)  | (\690(535)  | \689(1125) ),
  \2642(1304)  = ~\2467(1275) ,
  \2328(1101)  = \1912(1076)  & \2285(241) ,
  \630(246)  = \905(155)  & \540(65) ,
  \675(178)  = \802(100) ,
  \1992(966)  = ~\1967(882) ,
  \1640(1289)  = ~\1642(1259) ,
  \1978(933)  = \1975(790) ,
  \1401(776)  = \1393(666)  & \294(39) ,
  \2698(556)  = ~\870(443) ,
  \1608(1089)  = \1607(1033)  | \1606(1032) ,
  \691(524)  = \688(428)  & \540(65) ,
  \1012(386)  = \1009(318)  & \107(12) ,
  \3044(245)  = ~\3040(152) ,
  \1365(632)  = ~\1147(508) ,
  \2975(498)  = \557(366) ,
  \647(391)  = ~\3102(249)  | ~\3095(72) ,
  \3251(1208)  = ~\3245(1172) ,
  \3417(1431)  = ~\3411(1403) ,
  \3312(1290)  = ~\3308(1260) ,
  \3093(171)  = ~\3087(90) ,
  \2051(104)  = ~\33(3) ,
  \2046(1060)  = ~\2037(1003)  & ~\2034(1009) ,
  \3260(1436)  = ~\3256(1409) ,
  \1809(343)  = \1808(195)  & (\13(1)  & \1(0) ),
  \1716(294)  = ~\1681(192) ,
  \3313(1336)  = \2519(1300) ,
  \1287(817)  = \1279(707)  & \143(19) ,
  \2616(1421)  = ~\3410(1330)  | ~\3403(1402) ,
  \1743(496)  = \1742(364)  | (\1741(230)  | \1740(385) ),
  \2324(1202)  = ~\3138(1051)  | ~\3131(1184) ,
  \1328(614)  = ~\1111(506) ,
  \2990(481)  = ~\2986(355) ,
  \2674(1549)  = ~\2677(1514)  | ~\2676(1533) ,
  \2323(1238)  = ~\3137(1222)  | ~\3134(986) ,
  \1406(849)  = \1398(714)  & \517(70) ,
  \2314(1205)  = ~\2103(1110)  | (~\2210(1107)  | (~\2157(1169)  | ~\2257(1053) )),
  \1953(452)  = \1773(345)  & \1834(215) ,
  \2273(1218)  = ~\1993(1061)  | (~\1947(1170)  | ~\1895(1115) ),
  \2671(1550)  = ~\3449(1525)  | ~\3446(1495) ,
  \365(1570)  = \951(1564)  | (\947(910)  | \944(969) ),
  \1628(448)  = ~\1572(334) ,
  \2856(1690)  = ~\2855(1679)  | ~\2854(1685) ,
  \3303(1340)  = ~\3301(1306)  | ~\3298(1316) ,
  \1808(195)  = ~\788(109) ,
  \2895(1659)  = ~\3555(1646)  | ~\3552(1610) ,
  \2955(222)  = ~\2953(138)  | ~\2950(55) ,
  \2513(1343)  = \2426(1307)  & (\2433(1251)  & \2439(1281) ),
  \1480(607)  = ~\1186(505) ,
  \1589(306)  = ~\1512(193) ,
  \575(586)  = ~\2990(481)  | ~\2983(359) ,
  \1952(337)  = ~\1834(215) ,
  \1479(687)  = ~\1177(515) ,
  \1302(903)  = \1294(612)  & \432(99) ,
  \3137(1222)  = ~\3131(1184) ,
  \2887(1647)  = ~\3548(1621)  | ~\3541(1632) ,
  \905(155)  = \851(68)  & (\848(73)  & \842(77) ),
  \3435(1528)  = ~\2578(1511) ,
  \2312(1175)  = ~\2152(1149)  | ~\2103(1110) ,
  \2532(1303)  = ~\2467(1275)  | (~\2419(1288)  | ~\2409(1285) ),
  \1920(281)  = ~\807(181) ,
  \1563(329)  = ~\784(191)  | (~\732(117)  | ~\724(119) ),
  \1369(856)  = \1361(600)  & \504(76) ,
  \1274(659)  = ~\1075(512) ,
  \2811(1393)  = \2804(575)  & \1680(1359) ,
  \3127(1221)  = ~\3121(1183) ,
  \1583(1021)  = \1512(193)  & \1409(917) ,
  \1655(437)  = ~\1563(329) ,
  \1873(741)  = \1722(502)  & \1812(458) ,
  \3227(1210)  = ~\3221(1173) ,
  \2690(1611)  = \2687(1388)  | (\2684(1596)  | \2681(1574) ),
  \2706(1444)  = \2699(569)  & \1626(1417) ,
  \359(587)  = \923(482)  | (\920(361)  | \917(549) ),
  \1281(643)  = ~\1159(510) ,
  \1493(753)  = \1485(655)  & \322(43) ,
  \1588(1084)  = \1587(1023)  | \1586(1022) ,
  \914(440)  = ~\855(330) ,
  \600(1012)  = \597(960) ,
  \2664(1544)  = ~\3433(1529)  | ~\3430(1537) ,
  \2787(574)  = \870(443)  & \956(346) ,
  \1667(1280)  = ~\1669(1252) ,
  \3467(1591)  = \2780(1580) ,
  \2110(455)  = \1773(345)  & \1834(215) ,
  \2396(1253)  = ~\2395(1191)  | ~\2394(1228) ,
  \3539(1692)  = ~\3533(1687) ,
  \587(54)  = \264(35)  | \257(34) ,
  \3323(1138)  = \2458(1096) ,
  \1349(647)  = ~\1159(510) ,
  \1485(655)  = ~\1231(511) ,
  \3514(1634)  = ~\3510(1625) ,
  \2432(1189)  = ~\3228(1040)  | ~\3221(1173) ,
  \1761(352)  = \1758(300)  & \294(39) ,
  \1625(732)  = \1620(565)  & \456(94) ,
  \1653(1357)  = ~\1652(1090)  & (~\1650(1322)  & ~\1648(1131) ),
  \1260(610)  = ~\1111(506) ,
  \2957(53)  = \264(35) ,
  \1380(697)  = ~\1204(517) ,
  \3045(383)  = ~\3043(254)  | ~\3040(152) ,
  \2048(1111)  = \2047(1072)  & \2046(1060) ,
  \2184(747)  = \1764(488)  & \1794(460) ,
  \2687(1388)  = \2680(568)  & \1617(1356) ,
  \1963(881)  = \1960(540)  | (\1957(407)  | \1954(736) ),
  \1347(711)  = ~\1135(518) ,
  \3146(1167)  = ~\3142(1143) ,
  \2880(1620)  = \2690(1611)  & \2871(128) ,
  \2346(1256)  = ~\2345(1194)  | ~\2344(1231) ,
  \1367(799)  = \1359(664)  & \159(21) ,
  \3112(1464)  = ~\3268(1414)  | ~\3261(1438) ,
  \2512(1314)  = \2415(1287)  & \2495(1283) ,
  \1755(225)  = \1752(188)  & \244(32) ,
  \1258(674)  = ~\1087(514) ,
  \3069(1073)  = ~\3063(1013) ,
  \3082(165)  = \898(84) ,
  \1069(311)  = \1057(197)  & \1050(113) ,
  \2874(129)  = ~\2868(50)  & ~\2865(61) ,
  \2079(745)  = \1750(494)  & \1794(460) ,
  \1924(791)  = \1923(742)  | (\1922(478)  | \1921(495) ),
  \2827(1630)  = ~\3474(1618)  | ~\3467(1591) ,
  \678(275)  = ~\675(178) ,
  \1006(409)  = \1003(325)  & \833(86) ,
  \3379(1478)  = \2586(1459) ,
  \3369(1477)  = ~\3363(1458) ,
  \1409(917)  = ~\1408(783)  & (~\1407(839)  & (~\1406(849)  & (~\1405(858)  & (~\1404(868)  & (~\1403(878)  & (~\1402(889)  & ~\1401(776) )))))),
  \2966(220)  = ~\2964(131)  | ~\2957(53) ,
  \1030(1442)  = ~\938(722)  & (~\933(1419)  & ~\929(734) ),
  \2854(1685)  = ~\3523(1680)  | ~\3520(1661) ,
  \1307(954)  = ~\1306(821)  & (~\1305(816)  & (~\1304(810)  & (~\1303(803)  & (~\1302(903)  & (~\1301(893)  & (~\1300(883)  & ~\1299(825) )))))),
  \1418(769)  = \1410(667)  & \303(40) ,
  \1433(636)  = ~\1222(509) ,
  \917(549)  = \914(440)  & \650(273) ,
  \1060(243)  = \1054(196)  & \200(25) ,
  \717(120)  = \13(1) ,
  \1603(1031)  = \1512(193)  & \1494(912) ,
  \1356(906)  = \1348(631)  & \432(99) ,
  \369(1321)  = \[6] ,
  \2519(1300)  = \2518(1274)  | \2455(1095) ,
  \1487(844)  = \1479(687)  & \530(66) ,
  \1666(1133)  = \1663(583)  & \1604(1088) ,
  \3272(1262)  = ~\3130(1201)  | ~\3129(1237) ,
  \938(722)  = \928(576)  & \630(246) ,
  \1323(815)  = \1315(645)  & \143(19) ,
  \3071(1014)  = \591(965) ,
  \2202(994)  = \2193(923)  & (\2177(846)  & \190(24) ),
  \3498(1636)  = ~\3494(1627) ,
  \3366(1364)  = \2567(1333) ,
  \954(1532)  = ~\3119(1518)  | ~\3116(1494) ,
  \1600(1087)  = \1599(1029)  | \1598(1028) ,
  \3035(394)  = ~\3033(258)  | ~\3030(161) ,
  \2681(1574)  = \2678(462)  & \2549(1559) ,
  \2647(1372)  = ~\2645(1305)  & ~\2643(1328) ,
  \3147(1242)  = \2325(1204) ,
  \1342(663)  = ~\1075(512) ,
  \1662(1418)  = ~\1661(1126)  & (~\1659(1386)  & ~\1657(1132) ),
  \1437(860)  = \1429(604)  & \504(76) ,
  \1498(624)  = ~\1195(507) ,
  \1415(715)  = ~\1213(519) ,
  \3170(1045)  = ~\3166(980) ,
  \2734(558)  = ~\870(443) ,
  \2371(1199)  = ~\3204(1049)  | ~\3197(1177) ,
  \2236(748)  = \1771(485)  & \1794(460) ,
  \3465(1505)  = ~\3459(1485) ,
  \402(1718)  = \[21] ,
  \1883(1011)  = \1877(937)  & (\1862(899)  & \169(22) ),
  \460(89)  = \68(8) ,
  \1930(936)  = ~\1924(791) ,
  \1909(545)  = \1902(451)  & (\1829(214)  & \58(7) ),
  \2603(1488)  = ~\2602(1449)  | ~\2601(1471) ,
  \1255(833)  = \1247(641)  & \125(15) ,
  \1243(609)  = ~\1111(506) ,
  \617(536)  = \613(423)  & \501(79) ,
  \2536(1440)  = ~\3259(1383)  | ~\3256(1409) ,
  \1756(360)  = \1753(290)  & \250(33) ,
  \788(109)  = \41(4)  & \33(3) ,
  \3459(1485)  = \2814(1467) ,
  \3013(174)  = ~\3007(97) ,
  \1271(827)  = \1263(626)  & \132(17) ,
  \2716(464)  = ~\956(346) ,
  \1453(861)  = \1445(685)  & \504(76) ,
  \1623(1387)  = \1619(447)  & \1622(1351) ,
  \2931(60)  = \226(29) ,
  \897(168)  = ~\836(85)  | (~\831(92)  | ~\826(96) ),
  \1204(517)  = \1120(376) ,
  \911(724)  = ~\910(527) ,
  \2098(989)  = \2085(928)  & (\2072(863)  & \200(25) ),
  \2062(395)  = ~\1773(345)  & ~\87(10) ,
  \907(67)  = \107(12) ,
  \1530(302)  = ~\794(182)  | ~\776(107) ,
  \2844(1662)  = ~\2843(1651)  | ~\2842(1638) ,
  \2668(1576)  = ~\2667(1569) ,
  \2272(1182)  = ~\1942(1154)  | ~\1895(1115) ,
  \432(99)  = \50(6) ,
  \2298(237)  = \343(47)  & (\213(26)  & \2278(207) ),
  \2495(1283)  = \2491(1255) ,
  \3110(251)  = ~\3106(154) ,
  \501(79)  = ~\87(10) ,
  \3513(1613)  = ~\3507(1598) ,
  \1156(373)  = ~\1060(243)  | ~\1038(148) ,
  \1834(215)  = \1827(122)  & \1826(123) ,
  \932(1371)  = \2645(1305)  | \2643(1328) ,
  \1022(206)  = ~\741(116) ,
  \1618(578)  = ~\1545(470) ,
  \2970(491)  = \562(363) ,
  \3182(982)  = \2354(946) ,
  \3166(980)  = \2341(945) ,
  \981(314)  = ~\759(198) ,
  \2877(217)  = \2874(129) ,
  \2415(1287)  = \2359(1258) ,
  \2255(987)  = \2242(919)  & (\2229(836)  & \200(25) ),
  \2593(1489)  = ~\3386(1423)  | ~\3379(1478) ,
  \2623(1470)  = ~\2622(1422)  | ~\2621(1448) ,
  \2210(1107)  = \2209(1068)  & \2208(1056) ,
  \1439(841)  = \1431(700)  & \530(66) ,
  \586(356)  = ~\554(219)  | ~\553(227) ,
  \1405(858)  = \1397(698)  & \504(76) ,
  \1629(566)  = \1572(334)  & \1545(470) ,
  \3219(1267)  = ~\3213(1240) ,
  \1262(706)  = ~\1135(518) ,
  \1326(678)  = ~\1087(514) ,
  \1353(875)  = \1345(615)  & \483(81) ,
  \802(100)  = ~\45(5) ,
  \569(796)  = ~\2981(592)  | ~\2978(492) ,
  \3047(546)  = ~\3016(419)  | ~\3015(270) ,
  \3305(1380)  = ~\2535(1338)  | (~\2534(1335)  | ~\2533(1193) ),
  \1497(608)  = ~\1186(505) ,
  \2341(945)  = \1963(881)  & \2289(239) ,
  \408(1660)  = \2930(1649)  & \213(26) ,
  \649(723)  = \648(526)  & \530(66) ,
  \1455(842)  = \1447(621)  & \530(66) ,
  \2375(1097)  = \2120(1069)  & \2298(237) ,
  \1421(859)  = \1413(619)  & \504(76) ,
  \1764(488)  = \1763(358)  | (\1762(223)  | \1761(352) ),
  \1072(374)  = ~\1069(311)  | ~\1043(149) ,
  \1249(806)  = \1241(673)  & \159(21) ,
  \2963(133)  = ~\2957(53) ,
  \3531(1691)  = ~\3525(1686) ,
  \1250(813)  = \1242(593)  & \150(20) ,
  \668(425)  = \806(293)  & \804(303) ,
  \2358(1196)  = ~\3178(1046)  | ~\3171(1178) ,
  \2658(1575)  = ~\2638(1483)  & ~\2555(1566) ,
  \492(80)  = \87(10) ,
  \901(542)  = ~\904(412)  | ~\903(264) ,
  \1745(187)  = ~\1699(105) ,
  \3103(71)  = \97(11) ,
  \386(1602)  = ~\2765(1590) ,
  \2699(569)  = \870(443)  & \956(346) ,
  \2585(1411)  = ~\3312(1290)  | ~\3305(1380) ,
  \1471(843)  = \1463(606)  & \530(66) ,
  \1501(640)  = ~\1222(509) ,
  \1534(431)  = ~\1530(302) ,
  \2362(1234)  = ~\3185(1217)  | ~\3182(982) ,
  \1282(829)  = \1274(659)  & \128(16) ,
  \903(264)  = ~\3093(171)  | ~\3090(166) ,
  \1231(511)  = \1156(373) ,
  \1829(214)  = \1(0)  | \1828(110) ,
  \1856(417)  = ~\1773(345)  & ~\50(6) ,
  \2983(359)  = ~\2956(224)  | ~\2955(222) ,
  \2805(1446)  = \2802(469)  & \2626(1395) ,
  \2780(1580)  = \2777(1445)  | (\2774(1572)  | \2771(1523) ),
  \2670(1551)  = ~\3442(1519)  | ~\3435(1528) ,
  \2760(1391)  = \2753(572)  & \1653(1357) ,
  \1057(197)  = ~\1051(112) ,
  \2667(1569)  = ~\2670(1551)  | ~\2669(1563) ,
  \2757(1579)  = \2752(559)  & \2663(1567) ,
  \2150(1102)  = \2137(925)  & (\2124(1070)  & \200(25) ),
  \1322(809)  = \1314(629)  & \150(20) ,
  \2021(283)  = ~\807(181) ,
  \1488(778)  = \1480(607)  & \283(38) ,
  \799(101)  = \45(5) ,
  \3451(1487)  = ~\2623(1470) ,
  \3361(1476)  = ~\3355(1457) ,
  \1407(839)  = \1399(634)  & \530(66) ,
  \353(405)  = \[0] ,
  \1298(644)  = ~\1159(510) ,
  \2167(384)  = ~\1773(345)  & ~\107(12) ,
  \1397(698)  = ~\1204(517) ,
  \1410(667)  = ~\1168(513) ,
  \2718(570)  = \870(443)  & \956(346) ,
  \1277(611)  = ~\1111(506) ,
  \1826(123)  = ~\13(1)  | ~\1(0) ,
  \1108(371)  = ~\1066(312)  | ~\1038(148) ,
  \2004(737)  = \2002(338)  & \1000(538) ,
  \759(198)  = \20(2)  | \758(108) ,
  \2553(1531)  = ~\3346(1453)  | ~\3339(1517) ,
  \3302(1348)  = ~\3298(1316) ,
  \589(880)  = ~\3053(731)  | ~\3050(539) ,
  \2896(1648)  = ~\3556(1622)  | ~\3549(1633) ,
  \1582(1020)  = \1581(304)  & \1273(956) ,
  \3497(1554)  = ~\3491(1539) ,
  \2349(1232)  = ~\3169(1220)  | ~\3166(980) ,
  \2859(1708)  = ~\3539(1692)  | ~\3536(1698) ,
  \898(84)  = \68(8) ,
  \2313(1209)  = ~\2205(1055)  | (~\2157(1169)  | ~\2103(1110) ),
  \1656(552)  = \1563(329)  & \1554(471) ,
  \3130(1201)  = ~\3128(1050)  | ~\3121(1183) ,
  \3378(1299)  = ~\3374(1273) ,
  \3002(971)  = \579(939) ,
  \2739(1501)  = \2734(558)  & \2581(1472) ,
  \3520(1661)  = ~\3516(1650)  | ~\3515(1635) ,
  \855(330)  = ~\736(118)  | (~\721(211)  | ~\707(127) ),
  \1676(1282)  = ~\1678(1254) ,
  \1508(755)  = \1500(720)  & \317(42) ,
  \1542(348)  = ~\1541(151)  | (~\721(211)  | ~\707(127) ),
  \3134(986)  = \2320(948) ,
  \1734(232)  = \1731(185)  & \226(29) ,
  \1605(310)  = ~\1512(193) ,
  \1010(326)  = \759(198)  & \741(116) ,
  \2833(1681)  = ~\2832(1674)  | ~\2831(1664) ,
  \2445(1098)  = \2293(238)  & \1993(1061) ,
  \906(156)  = ~\851(68)  | (~\848(73)  | ~\842(77) ),
  \1423(840)  = \1415(715)  & \530(66) ,
  \1382(633)  = ~\1222(509) ,
  \591(965)  = ~\590(891)  | ~\589(880) ,
  \3053(731)  = ~\3047(546) ,
  \2511(1313)  = \2409(1285)  & (\2419(1288)  & \2495(1283) ),
  \2455(1095)  = \2302(236)  & \2205(1055) ,
  \2697(463)  = ~\956(346) ,
  \2531(1312)  = ~\2451(1142)  | ~\2409(1285) ,
  \2131(746)  = \1757(490)  & \1794(460) ,
  \1622(1351)  = ~\1624(1318) ,
  \2483(999)  = \2478(64)  & (\2477(921)  & (\2476(924)  & (\2475(927)  & \2474(930) ))),
  \1288(822)  = \1280(627)  & \137(18) ,
  \2660(1584)  = \2659(1568)  | \2658(1575) ,
  \2592(1508)  = ~\3385(1496)  | ~\3382(1396) ,
  \2797(1582)  = \2794(1392)  | (\2791(1573)  | \2788(1503) ),
  \2007(401)  = ~\1773(345)  & ~\77(9) ,
  \2956(224)  = ~\2954(135)  | ~\2947(56) ,
  \3528(1697)  = \2856(1690) ,
  \2040(996)  = \2031(932)  & (\2017(872)  & \190(24) ),
  \1359(664)  = ~\1075(512) ,
  \2526(1370)  = ~\2467(1275)  | (~\2419(1288)  | (~\2406(1284)  | ~\2401(1350) )),
  \595(837)  = ~\3061(725)  | ~\3058(522) ,
  \603(1120)  = ~\3077(1074)  | ~\3074(1067) ,
  \1735(365)  = \1732(287)  & \232(30) ,
  \1001(203)  = ~\741(116) ,
  \1345(615)  = ~\1111(506) ,
  \608(1185)  = ~\607(1158)  | ~\606(1118) ,
  \707(127)  = \1(0) ,
  \3568(1694)  = \2913(1688) ,
  \3102(249)  = ~\3098(153) ,
  \2177(846)  = ~\2170(525)  & (~\2167(384)  & ~\2164(739) ),
  \2288(240)  = ~\213(26)  | ~\2278(207) ,
  \1029(588)  = ~\923(482)  & (~\920(361)  & ~\917(549) ),
  \2190(922)  = \2185(786) ,
  \980(200)  = ~\741(116) ,
  \2219(380)  = ~\1773(345)  & ~\116(13) ,
  \375(1624)  = \2690(1611) ,
  \1496(688)  = ~\1177(515) ,
  \1974(743)  = \1736(500)  & \1812(458) ,
  \1599(1029)  = \1512(193)  & \1477(913) ,
  \3211(1266)  = ~\3205(1239) ,
  \2579(1450)  = ~\3377(1433)  | ~\3374(1273) ,
  \2612(1272)  = \2396(1253)  & \330(46) ,
  \3386(1423)  = ~\3382(1396) ,
  \1889(998)  = \1880(938)  & (\1866(900)  & \190(24) ),
  \1744(298)  = ~\1681(192) ,
  \1895(1115)  = \1894(1078)  & \1893(1064) ,
  \1472(779)  = \1464(622)  & \283(38) ,
  \2156(1145)  = \2151(1122)  | (\2150(1102)  | \2149(1104) ),
  \1675(1134)  = \1672(584)  & \1608(1089) ,
  \1602(1030)  = \1601(309)  & \1358(951) ,
  \2099(963)  = ~\2072(863) ,
  \2937(146)  = ~\2931(60) ,
  \1772(212)  = ~\731(121) ,
  \2615(1447)  = ~\3409(1430)  | ~\3406(1297) ,
  \701(523)  = \696(429)  & \634(247) ,
  \384(1553)  = \[10] ,
  \483(81)  = \77(9) ,
  \1645(581)  = ~\1554(471) ,
  \1456(780)  = \1448(701)  & \283(38) ,
  \1016(319)  = ~\759(198) ,
  \3040(152)  = \540(65) ,
  \645(890)  = \644(269)  | \641(728) ,
  \2925(1629)  = \2694(1612)  & (\2713(1588)  & (\2730(1600)  & \2748(1522) )),
  \2950(55)  = \257(34) ,
  \2293(238)  = ~\343(47)  | (~\213(26)  | ~\2278(207) ),
  \1732(287)  = \1699(105)  & \1681(192) ,
  \3422(1311)  = \2439(1281) ,
  \1615(1263)  = ~\2324(1202)  | ~\2323(1238) ,
  \1366(648)  = ~\1159(510) ,
  \663(1124)  = ~\662(550)  & ~\661(1080) ,
  \3058(522)  = ~\3046(387)  | ~\3045(383) ,
  \3236(1041)  = ~\3232(976) ,
  \1679(1188)  = \1674(554)  & \692(1157) ,
  \3245(1172)  = \2388(1147) ,
  \2572(1510)  = ~\2571(1473)  | ~\2570(1491) ,
  \550(136)  = ~\504(76)  | ~\257(34) ,
  \545(147)  = ~\432(99)  | ~\226(29) ,
  \2205(1055)  = \2199(1001)  | \2196(1007) ,
  \1740(385)  = \1737(297)  & \107(12) ,
  \2728(1599)  = \2725(1389)  | (\2722(1586)  | \2719(1538) ),
  \401(1716)  = ~\2860(1710)  | ~\2859(1708) ,
  \986(958)  = \985(378)  | (\984(408)  | \983(908) ),
  \1438(851)  = \1430(620)  & \517(70) ,
  \1256(957)  = ~\1255(833)  & (~\1254(831)  & (~\1253(828)  & (~\1252(824)  & (~\1251(819)  & (~\1250(813)  & (~\1249(806)  & ~\1248(834) )))))),
  \1871(499)  = \1870(280)  & (\226(29)  & \1817(459) ),
  \1364(712)  = ~\1135(518) ,
  \3046(387)  = ~\3044(245)  | ~\3037(157) ,
  \1291(660)  = ~\1075(512) ,
  \3043(254)  = ~\3037(157) ,
  \1299(825)  = \1291(660)  & \132(17) ,
  \2672(1524)  = ~\3450(1515)  | ~\3443(1507) ,
  \1019(382)  = \1016(319)  & \116(13) ,
  \2544(1400)  = \2508(1381)  & \330(46) ,
  \1279(707)  = ~\1135(518) ,
  \2939(58)  = \238(31) ,
  \1435(763)  = \1427(668)  & \311(41) ,
  \3304(1373)  = ~\3302(1348)  | ~\3295(1276) ,
  \1760(291)  = \1699(105)  & \1681(192) ,
  \2351(1152)  = \2048(1111) ,
  \3155(1180)  = \2338(1153) ,
  \3517(1672)  = \2844(1662) ,
  \1454(852)  = \1446(605)  & \517(70) ,
  \848(73)  = ~\97(11) ,
  \1400(650)  = ~\1231(511) ,
  \1942(1154)  = \1936(1113)  | \1933(1117) ,
  \2320(948)  = \1862(899)  & \2285(241) ,
  \1275(675)  = ~\1087(514) ,
  \3142(1143)  = \2328(1101) ,
  \1724(184)  = ~\1699(105) ,
  \3111(1482)  = ~\3267(1460)  | ~\3264(1384) ,
  \1408(783)  = \1400(650)  & \283(38) ,
  \597(960)  = ~\596(854)  | ~\595(837) ,
  \3186(1047)  = ~\3182(982) ,
  \1817(459)  = ~\1809(343) ,
  \1339(801)  = \1331(630)  & \159(21) ,
  \1470(853)  = \1462(686)  & \517(70) ,
  \2085(928)  = \2080(788) ,
  \2350(1195)  = ~\3170(1045)  | ~\3163(1181) ,
  \904(412)  = ~\3094(265)  | ~\3087(90) ,
  \1032(115)  = ~\20(2) ,
  \588(137)  = \587(54)  & \250(33) ,
  \1301(893)  = \1293(596)  & \447(95) ,
  \3185(1217)  = ~\3179(1179) ,
  \1554(471)  = \1542(348) ,
  \1659(1386)  = \1655(437)  & \1658(1342) ,
  \1758(300)  = ~\1681(192) ,
  \1450(637)  = ~\1222(509) ,
  \571(942)  = ~\570(798)  | ~\569(796) ,
  \3401(1454)  = ~\3395(1429) ,
  \1426(916)  = ~\1425(775)  & (~\1424(782)  & (~\1423(840)  & (~\1422(850)  & (~\1421(859)  & (~\1420(869)  & (~\1419(879)  & ~\1418(769) )))))),
  \982(322)  = \759(198)  & \741(116) ,
  \3086(263)  = ~\3082(165) ,
  \3224(975)  = \2383(943) ,
  \2953(138)  = ~\2947(56) ,
  \1997(1075)  = \1992(966)  | (\1991(991)  | \1990(997) ),
  \357(1136)  = ~\583(1094)  | ~\582(1092) ,
  \2302(236)  = ~\343(47)  | (~\213(26)  | ~\2278(207) ),
  \1424(782)  = \1416(635)  & \283(38) ,
  \1324(953)  = ~\1323(815)  & (~\1322(809)  & (~\1321(802)  & (~\1320(904)  & (~\1319(894)  & (~\1318(884)  & (~\1317(873)  & ~\1316(820) )))))),
  \3552(1610)  = \2883(1595) ,
  \1933(1117)  = \1927(935)  & (\1912(1076)  & \169(22) ),
  \1614(1325)  = \1610(446)  & \1613(1293) ,
  \2973(591)  = ~\2967(497) ,
  \2625(1360)  = ~\3426(1344)  | ~\3419(51) ,
  \1020(398)  = \1017(327)  & \839(78) ,
  \3338(1452)  = ~\3334(1426) ,
  \2256(959)  = ~\2229(836) ,
  \1736(500)  = \1735(365)  | (\1734(232)  | \1733(389) ),
  \942(441)  = ~\855(330) ,
  \2400(1192)  = ~\3252(1043)  | ~\3245(1172) ,
  \2338(1153)  = \1998(1112) ,
  \1413(619)  = ~\1195(507) ,
  \2426(1307)  = ~\2425(1249)  | ~\2424(1277) ,
  \928(576)  = \893(216)  & \887(444) ,
  \2399(1229)  = ~\3251(1208)  | ~\3248(978) ,
  \991(404)  = \988(315)  & \77(9) ,
  \1427(668)  = ~\1168(513) ,
  \352(260)  = ~\625(167)  | ~\479(82) ,
  \2826(1617)  = ~\3473(1604)  | ~\3470(1601) ,
  \1527(284)  = ~\794(182)  | ~\784(191) ,
  \807(181)  = \798(102)  & \714(124) ,
  \2229(836)  = ~\2222(520)  & (~\2219(380)  & ~\2216(740) ),
  \1853(735)  = \1851(335)  & \979(543) ,
  \993(544)  = \992(418)  | (\991(404)  | \990(267) ),
  \3138(1051)  = ~\3134(986) ,
  \3470(1601)  = \2763(1589) ,
  \2843(1651)  = ~\3498(1636)  | ~\3491(1539) ,
  \1440(781)  = \1432(716)  & \283(38) ,
  \2137(925)  = \2132(787) ,
  \3128(1050)  = ~\3124(985) ,
  \3285(1413)  = ~\3283(1376)  | ~\3280(1349) ,
  \1672(584)  = ~\1554(471) ,
  \3286(1407)  = ~\3284(1382)  | ~\3277(1345) ,
  \2662(1548)  = \2650(1404)  & (\2594(1526)  & (\2603(1488)  & \2617(1469) )),
  \3560(1693)  = \2913(1688) ,
  \2626(1395)  = ~\2625(1360)  | ~\2624(1329) ,
  \1284(902)  = \1276(595)  & \432(99) ,
  \2401(1350)  = \2333(1317) ,
  \2424(1277)  = ~\3211(1266)  | ~\3208(1139) ,
  \3256(1409)  = \2508(1381) ,
  \1195(507)  = \1108(371) ,
  \1768(351)  = \1765(301)  & \303(40) ,
  \673(1082)  = \672(533)  | (\671(426)  | \669(1019) ),
  \1596(1086)  = \1595(1027)  | \1594(1026) ,
  \3079(91)  = \58(7) ,
  \2719(1538)  = \2716(464)  & \2572(1510) ,
  \823(180)  = \799(101)  & \704(126) ,
  \2387(1190)  = ~\3236(1041)  | ~\3229(1174) ,
  \442(98)  = ~\50(6) ,
  \2733(465)  = ~\956(346) ,
  \1535(422)  = \1530(302)  & \1527(284) ,
  \2853(1652)  = ~\3506(1637)  | ~\3499(1540) ,
  \3240(977)  = \2391(944) ,
  \3502(1628)  = \2839(1614) ,
  \3433(1529)  = ~\3427(1512) ,
  \3235(1211)  = ~\3229(1174) ,
  \1422(850)  = \1414(699)  & \517(70) ,
  \3124(985)  = \2320(948) ,
  \3154(1168)  = ~\3150(1144) ,
  \1399(634)  = ~\1222(509) ,
  \685(427)  = ~\806(293) ,
  \1412(603)  = ~\1186(505) ,
  \1922(478)  = \807(181)  & (\274(37)  & \1817(459) ),
  \1272(830)  = \1264(642)  & \128(16) ,
  \2474(930)  = ~\2080(788) ,
  \2539(1480)  = ~\3275(1461)  | ~\3272(1262) ,
  \2022(489)  = \2021(283)  & (\244(32)  & \1817(459) ),
  \2242(919)  = \2237(785) ,
  \831(92)  = ~\58(7) ,
  \2599(1527)  = ~\2598(1490)  | ~\2597(1509) ,
  \1300(883)  = \1292(676)  & \467(87) ,
  \2372(1203)  = \2157(1169) ,
  \2607(1301)  = ~\3329(1162)  | ~\3326(1279) ,
  \1591(1025)  = \1512(193)  & \1443(915) ,
  \1159(510)  = \1156(373) ,
  \1386(888)  = \1378(601)  & \467(87) ,
  \1370(866)  = \1362(616)  & \492(80) ,
  \2552(1546)  = ~\3345(1535)  | ~\3342(1427) ,
  \2666(1565)  = ~\2665(1558)  | ~\2664(1544) ,
  \2031(932)  = ~\2025(789) ,
  \1432(716)  = ~\1213(519) ,
  \956(346)  = \896(176)  & \890(125) ,
  \1489(771)  = \1481(623)  & \294(39) ,
  \3398(1332)  = \2514(1309)  & \330(46) ,
  \1671(1358)  = ~\1670(1225)  & (~\1668(1323)  & ~\1666(1133) ),
  \607(1158)  = ~\3070(1119)  | ~\3063(1013) ,
  \2725(1389)  = \2718(570)  & \1635(1355) ,
  \700(1160)  = \694(435)  & \663(1124) ,
  \1355(896)  = \1347(711)  & \447(95) ,
  \1670(1225)  = \1665(553)  & \703(1187) ,
  \2803(562)  = ~\870(443) ,
  \407(1657)  = \[18] ,
  \1343(679)  = ~\1087(514) ,
  \553(227)  = \548(141)  & (\547(143)  & (\546(145)  & \545(147) )),
  \1021(529)  = \1020(398)  | (\1019(382)  | \1018(253) ),
  \2478(64)  = \179(23) ,
  \2999(974)  = \571(942) ,
  \1048(62)  = ~\200(25) ,
  \1075(512)  = \1072(374) ,
  \1619(447)  = ~\1572(334) ,
  \2634(1416)  = \2629(1385)  & \2501(1353) ,
  \3264(1384)  = \2501(1353) ,
  \3284(1382)  = ~\3280(1349) ,
  \1624(1318)  = ~\2337(1265)  | ~\2336(1295) ,
  \2964(131)  = ~\2960(52) ,
  \2114(388)  = ~\1773(345)  & ~\97(11) ,
  \1147(508)  = \1144(372) ,
  \3516(1650)  = ~\3514(1634)  | ~\3507(1598) ,
  \1585(305)  = ~\1512(193) ,
  \3458(1455)  = ~\3454(1432) ,
  \2788(1503)  = \2785(468)  & \2617(1469) ,
  \1726(396)  = \1723(295)  & \87(10) ,
  \3077(1074)  = ~\3071(1014) ,
  \2584(1437)  = ~\3311(1408)  | ~\3308(1260) ,
  \1723(295)  = ~\1681(192) ,
  \1870(280)  = ~\807(181) ,
  \839(78)  = \87(10) ,
  \3308(1260)  = ~\3196(1198)  | ~\3195(1235) ,
  \3006(1037)  = ~\3002(971) ,
  \1312(693)  = ~\1123(516) ,
  \3395(1429)  = ~\3322(1401)  | ~\3321(1406) ,
  \3482(1665)  = ~\3478(1653) ,
  \951(1564)  = \943(445)  & \950(1547) ,
  \3387(1479)  = \2586(1459) ,
  \1431(700)  = ~\1204(517) ,
  \2517(1302)  = \2415(1287)  & \2467(1275) ,
  \3557(1695)  = \2910(1689) ,
  \3298(1316)  = \2415(1287) ,
  \2500(1319)  = \2268(1245)  & \2467(1275) ,
  \2146(1108)  = \2140(926)  & (\2120(1069)  & \179(23) ),
  \983(908)  = \980(200)  & \902(729) ,
  \1294(612)  = ~\1111(506) ,
  \1791(344)  = \1790(194)  & (\13(1)  & \1(0) ),
  \1827(122)  = ~\33(3)  | (~\20(2)  | ~\1(0) ),
  \1251(819)  = \1243(609)  & \143(19) ,
  \3195(1235)  = ~\3193(1212)  | ~\3190(983) ,
  \2832(1674)  = ~\3482(1665)  | ~\3475(1641) ,
  \1541(151)  = \169(22)  | \1540(111) ,
  \2431(1226)  = ~\3227(1210)  | ~\3224(975) ,
  \2525(1377)  = ~\2451(1142)  | (~\2406(1284)  | ~\2401(1350) ),
  \1598(1028)  = \1597(308)  & \1341(952) ,
  \2010(537)  = \2003(453)  & (\1829(214)  & \77(9) ),
  \3418(1331)  = ~\3414(1298) ,
  \2309(1206)  = \2262(1106)  & (\2210(1107)  & (\2157(1169)  & \2103(1110) )),
  \1646(436)  = ~\1563(329) ,
  \696(429)  = ~\806(293) ,
  \2523(1200)  = ~\2444(1166) ,
  \2608(1339)  = ~\3330(1310)  | ~\3323(1138) ,
  \2216(740)  = \2214(342)  & \1028(521) ,
  \3116(1494)  = \2538(1481)  & \330(46) ,
  \610(432)  = ~\804(303) ,
  \583(1094)  = ~\3006(1037)  | ~\2999(974) ,
  \702(530)  = \699(430)  & \526(69) ,
  \1750(494)  = \1749(362)  | (\1748(228)  | \1747(381) ),
  \2735(571)  = \870(443)  & \956(346) ,
  \392(1594)  = ~\2799(1583) ,
  \1509(752)  = \1501(640)  & \322(43) ,
  \1084(375)  = ~\1066(312)  | ~\1043(149) ,
  \400(1715)  = ~\2864(1709)  | ~\2863(1707) ,
  \2892(1678)  = ~\2891(1669) ,
  \2564(1435)  = ~\2563(1378)  | ~\2562(1410) ,
  \1643(727)  = \1638(567)  & \479(82) ,
  \2041(990)  = \2028(931)  & (\2017(872)  & \200(25) ),
  \3354(1365)  = ~\3350(1334) ,
  \1790(194)  = ~\788(109) ,
  \1616(733)  = \1611(564)  & \442(98) ,
  \2164(739)  = \2162(341)  & \1021(529) ,
  \1035(63)  = \190(24) ,
  \1417(651)  = ~\1231(511) ,
  \1457(773)  = \1449(717)  & \294(39) ,
  \3267(1460)  = ~\3261(1438) ,
  \2091(1008)  = \2085(928)  & (\2068(862)  & \169(22) ),
  \1812(458)  = \1809(343) ,
  \530(66)  = \116(13) ,
  \1996(1062)  = ~\1987(1004)  & ~\1984(1010) ,
  \1354(886)  = \1346(695)  & \467(87) ,
  \3549(1633)  = \2880(1620) ,
  \3443(1507)  = \2603(1488) ,
  \2518(1274)  = \2461(1137)  & \2433(1251) ,
  \929(734)  = \926(563)  & \650(273) ,
  \3205(1239)  = \2372(1203) ,
  \1473(772)  = \1465(702)  & \294(39) ,
  \1763(358)  = \1760(291)  & \257(34) ,
  \988(315)  = ~\759(198) ,
  \3030(161)  = \513(75) ,
  \990(267)  = \987(201)  & \836(85) ,
  \1467(638)  = ~\1222(509) ,
  \1049(114)  = \200(25)  & \20(2) ,
  \2157(1169)  = \2156(1145)  & \2155(1150) ,
  \2059(738)  = \2057(339)  & \1007(528) ,
  \2571(1473)  = ~\3362(1398)  | ~\3355(1457) ,
  \2581(1472)  = ~\2580(1425)  | ~\2579(1450) ,
  \1411(683)  = ~\1177(515) ,
  \2601(1471)  = ~\3401(1454)  | ~\3398(1332) ,
  \361(940)  = \[2] ,
  \3033(258)  = ~\3027(162) ,
  \916(442)  = \861(209)  & \855(330) ,
  \1320(904)  = \1312(693)  & \432(99) ,
  \2181(277)  = ~\816(179) ,
  \570(798)  = ~\2982(590)  | ~\2975(498) ,
  \1874(792)  = \1873(741)  | (\1872(479)  | \1871(499) ),
  \1500(720)  = ~\1213(519) ,
  \1762(223)  = \1759(189)  & \250(33) ,
  \1013(403)  = \1010(326)  & \77(9) ,
  \944(969)  = \941(333)  & \645(890) ,
  \1317(873)  = \1309(677)  & \483(81) ,
  \2370(1236)  = ~\3203(1213)  | ~\3200(984) ,
  \1350(807)  = \1342(663)  & \150(20) ,
  \1376(665)  = ~\1168(513) ,
  \2268(1245)  = \2265(1215) ,
  \3109(159)  = ~\3103(71) ,
  \2849(1673)  = ~\2848(1663) ,
  \1859(547)  = \1852(450)  & (\1829(214)  & \50(6) ),
  \1289(826)  = \1281(643)  & \132(17) ,
  \2530(1141)  = ~\2445(1098) ,
  \3489(1656)  = ~\3483(1642) ,
  \2960(52)  = \270(36) ,
  \2475(927)  = ~\2132(787) ,
  \2920(1711)  = ~\3563(1702)  | ~\3560(1693) ,
  \2638(1483)  = \2635(1465) ,
  \1673(439)  = ~\1563(329) ,
  \3095(72)  = \97(11) ,
  \2076(279)  = ~\823(180) ,
  \1043(149)  = ~\1035(63)  & ~\1032(115) ,
  \1916(1077)  = ~\1909(545)  & (~\1906(411)  & ~\1903(1034) ),
  \689(1125)  = \683(434)  & \681(1081) ,
  \1425(775)  = \1417(651)  & \294(39) ,
  \2124(1070)  = ~\2117(531)  & (~\2114(388)  & ~\2111(1035) ),
  \672(533)  = \668(425)  & \513(75) ,
  \2633(1420)  = \2632(1415)  & (\2505(1320)  & \330(46) ),
  \2938(144)  = ~\2934(59) ,
  \1880(938)  = ~\1874(792) ,
  \864(210)  = ~\724(119)  | ~\707(127) ,
  \867(332)  = ~\794(182)  | (~\736(118)  | (~\724(119)  | ~\707(127) )),
  \389(1592)  = ~\2782(1581) ,
  \902(729)  = ~\901(542) ,
  \1246(625)  = ~\1147(508) ,
  \1429(604)  = ~\1186(505) ,
  \3350(1334)  = \2511(1313)  & \330(46) ,
  \3454(1432)  = \2650(1404) ,
  \395(1486)  = ~\2816(1468) ,
  \2578(1511)  = ~\2577(1474)  | ~\2576(1492) ,
  \721(211)  = \717(120) ,
  \1362(616)  = ~\1111(506) ,
  \2170(525)  = \2163(456)  & (\2052(213)  & \107(12) ),
  \2111(1035)  = \2109(340)  & \1014(962) ,
  \3499(1540)  = \2745(1521) ,
  \3119(1518)  = ~\3113(1499) ,
  \1383(649)  = ~\1231(511) ,
  \1441(774)  = \1433(636)  & \294(39) ,
  \640(541)  = ~\643(413)  | ~\642(262) ,
  \724(119)  = ~\13(1) ,
  \2025(789)  = \2024(744)  | (\2023(476)  | \2022(489) ),
  \1443(915)  = ~\1442(768)  & (~\1441(774)  & (~\1440(781)  & (~\1439(841)  & (~\1438(851)  & (~\1437(860)  & (~\1436(870)  & ~\1435(763) )))))),
  \3253(1352)  = \2505(1320) ,
  \1452(758)  = \1444(669)  & \317(42) ,
  \2233(278)  = ~\816(179) ,
  \680(420)  = \675(178)  & \650(273) ,
  \1449(717)  = ~\1213(519) ,
  \1609(577)  = ~\1545(470) ,
  \2317(1156)  = \1895(1115) ,
  \1273(956)  = ~\1272(830)  & (~\1271(827)  & (~\1270(823)  & (~\1269(818)  & (~\1268(812)  & (~\1267(805)  & (~\1266(901)  & ~\1265(832) )))))),
  \1381(713)  = ~\1213(519) ,
  \2913(1688)  = ~\2838(1682) ,
  \642(262)  = ~\3085(172)  | ~\3082(165) ,
  \2017(872)  = ~\2010(537)  & (~\2007(401)  & ~\2004(737) ),
  \2289(239)  = \343(47)  & (\213(26)  & \2278(207) ),
  \3410(1330)  = ~\3406(1297) ,
  \356(1135)  = ~\620(1093)  | ~\619(1091) ,
  \1972(493)  = \1971(282)  & (\238(31)  & \1817(459) ),
  \1268(812)  = \1260(610)  & \150(20) ,
  \1005(392)  = \1002(317)  & \845(74) ,
  \2994(970)  = \579(939) ,
  \3301(1306)  = ~\3295(1276) ,
  \1017(327)  = \759(198)  & \741(116) ,
  \1242(593)  = ~\1099(504) ,
  \1296(708)  = ~\1135(518) ,
  \1038(148)  = \1035(63)  | \1032(115) ,
  \2538(1481)  = ~\2537(1463)  | ~\2536(1440) ,
  \551(134)  = ~\517(70)  | ~\264(35) ,
  \3276(1292)  = ~\3272(1262) ,
  \2541(1498)  = ~\2540(1462)  | ~\2539(1480) ,
  \826(96)  = ~\50(6) ,
  \546(145)  = ~\447(95)  | ~\232(30) ,
  \1954(736)  = \1952(337)  & \993(544) ,
  \1590(1024)  = \1589(306)  & \1307(954) ,
  \565(795)  = ~\2973(591)  | ~\2970(491) ,
  \3290(1315)  = \2409(1285) ,
  \3446(1495)  = \2647(1372)  & \2617(1469) ,
  \1014(962)  = \1013(403)  | (\1012(386)  | \1011(909) ),
  \943(445)  = \855(330)  & \864(210) ,
  \1384(784)  = \1376(665)  & \283(38) ,
  \3362(1398)  = ~\3358(1363) ,
  \3382(1396)  = \2589(1362) ,
  \3208(1139)  = \2375(1097) ,
  \1361(600)  = ~\1099(504) ,
  \1329(694)  = ~\1123(516) ,
  \3466(1606)  = ~\3462(1593) ,
  \1000(538)  = \999(415)  | (\998(397)  | \997(259) ),
  \2675(1562)  = ~\2674(1549) ,
  \2490(1230)  = \2485(369)  & \2309(1206) ,
  \2203(988)  = \2190(922)  & (\2177(846)  & \200(25) ),
  \2391(944)  = \2225(835)  & \2298(237) ,
  \362(1441)  = \938(722)  | (\933(1419)  | \929(734) ),
  \1374(907)  = \1366(648)  & \432(99) ,
  \1008(204)  = ~\741(116) ,
  \2128(276)  = ~\816(179) ,
  \2555(1566)  = ~\2554(1560) ,
  \3280(1349)  = \2333(1317) ,
  \1680(1359)  = ~\1679(1188)  & (~\1677(1324)  & ~\1675(1134) ),
  \860(208)  = \736(118)  & (\724(119)  & \707(127) ),
  \1448(701)  = ~\1204(517) ,
  \3541(1632)  = \2880(1620) ,
  \2954(135)  = ~\2950(55) ,
  \2484(1052)  = \2483(999)  | \2482(949) ,
  \1341(952)  = ~\1340(808)  & (~\1339(801)  & (~\1338(905)  & (~\1337(895)  & (~\1336(885)  & (~\1335(874)  & (~\1334(864)  & ~\1333(814) )))))),
  \3449(1525)  = ~\3443(1507) ,
  \2043(1059)  = \2037(1003)  | \2034(1009) ,
  \2665(1558)  = ~\3434(1552)  | ~\3427(1512) ,
  \2540(1462)  = ~\3276(1292)  | ~\3269(1439) ,
  \845(74)  = \97(11) ,
  \3330(1310)  = ~\3326(1279) ,
  \2567(1333)  = \2512(1314)  & \330(46) ,
  \1292(676)  = ~\1087(514) ,
  \2524(1375)  = ~\2445(1098)  | ~\2401(1350) ,
  \1537(1018)  = \1534(431)  & \1392(918) ,
  \616(424)  = ~\806(293) ,
  \1752(188)  = ~\1699(105) ,
  \2357(1233)  = ~\3177(1216)  | ~\3174(981) ,
  \987(201)  = ~\741(116) ,
  \1387(877)  = \1379(617)  & \483(81) ,
  \1444(669)  = ~\1168(513) ,
  \2752(559)  = ~\870(443) ,
  \2222(520)  = \2215(457)  & (\2052(213)  & \116(13) ),
  \3442(1519)  = ~\3438(1500) ,
  \1026(354)  = \1023(320)  & \283(38) ,
  \3005(1039)  = ~\2999(974) ,
  \1886(1005)  = \1880(938)  & (\1862(899)  & \179(23) ),
  \567(941)  = ~\566(797)  | ~\565(795) ,
  \3283(1376)  = ~\3277(1345) ,
  \3536(1698)  = \2856(1690) ,
  \1739(288)  = \1699(105)  & \1681(192) ,
  \3475(1641)  = \2823(1631) ,
  \1120(376)  = ~\1063(242)  | ~\1043(149) ,
  \2173(845)  = \2170(525)  | (\2167(384)  | \2164(739) ),
  \2679(555)  = ~\870(443) ,
  \3548(1621)  = ~\3544(1609) ,
  \2548(1530)  = ~\3338(1452)  | ~\3331(1516) ,
  \2433(1251)  = ~\2432(1189)  | ~\2431(1226) ,
  \2182(483)  = \2181(277)  & (\264(35)  & \1799(461) ),
  \1990(997)  = \1981(934)  & (\1967(882)  & \190(24) ),
  \2694(1612)  = ~\2687(1388)  & (~\2684(1596)  & ~\2681(1574) ),
  \3394(1424)  = ~\3390(1397) ,
  \1828(110)  = ~\20(2) ,
  \3293(1379)  = ~\3287(1346) ,
  \3066(1066)  = \600(1012) ,
  \2771(1523)  = \2768(467)  & \2603(1488) ,
  \1747(381)  = \1744(298)  & \116(13) ,
  \1018(253)  = \1015(205)  & \851(68) ,
  \1719(402)  = \1716(294)  & \77(9) ,
  \576(793)  = ~\575(586)  | ~\574(585) ,
  \2278(207)  = \732(117)  & (\717(120)  & \704(126) ),
  \1647(551)  = \1563(329)  & \1554(471) ,
  \1267(805)  = \1259(594)  & \159(21) ,
  \1430(620)  = ~\1195(507) ,
  \1261(690)  = ~\1123(516) ,
  \3441(1543)  = ~\3435(1528) ,
  \3334(1426)  = \2544(1400) ,
  \2485(369)  = \2293(238) ,
  \998(397)  = \995(316)  & \839(78) ,
  \3339(1517)  = \2541(1498) ,
  \1314(629)  = ~\1147(508) ,
  \3054(726)  = ~\3050(539) ,
  \2558(1493)  = ~\2557(1451)  | ~\2556(1475) ,
  \1771(485)  = \1770(357)  | (\1769(221)  | \1768(351) ),
  \2967(497)  = \557(366) ,
  \2598(1490)  = ~\3394(1424)  | ~\3387(1479) ,
  \1538(548)  = \1535(422)  & \442(98) ,
  \2557(1451)  = ~\3354(1365)  | ~\3347(1434) ,
  \582(1092)  = ~\3005(1039)  | ~\3002(971) ,
  \372(1243)  = \[5] ,
  \2921(1701)  = ~\3564(1699)  | ~\3557(1695) ,
  \1890(992)  = \1877(937)  & (\1866(900)  & \200(25) ),
  \1428(684)  = ~\1177(515) ,
  \1511(911)  = ~\1510(750)  & (~\1509(752)  & (~\1508(755)  & (~\1507(759)  & (~\1506(764)  & (~\1505(770)  & (~\1504(777)  & ~\1503(749) )))))),
  \3406(1297)  = \2612(1272) ,
  \3244(1042)  = ~\3240(977) ,
  \2802(469)  = ~\956(346) ,
  \1587(1023)  = \1512(193)  & \1426(916) ,
  \1927(935)  = \1924(791) ,
  \2103(1110)  = \2102(1071)  & \2101(1058) ,
  \2617(1469)  = ~\2616(1421)  | ~\2615(1447) ,
  \1741(230)  = \1738(186)  & \232(30) ,
  \2838(1682)  = ~\2837(1675)  | ~\2836(1666) ,
  \2748(1522)  = ~\2742(1390)  & (~\2739(1501)  & ~\2736(1502) ),
  \1504(777)  = \1496(688)  & \283(38) ,
  \1894(1078)  = \1891(967)  | (\1890(992)  | \1889(998) ),
  \758(108)  = ~\33(3) ,
  \3481(1655)  = ~\3475(1641) ,
  \870(443)  = \867(332) ,
  \2052(213)  = \1(0)  | \2051(104) ,
  \3204(1049)  = ~\3200(984) ,
  \3287(1346)  = \2517(1302)  | \2448(1099) ,
  \2537(1463)  = ~\3260(1436)  | ~\3253(1352) ,
  \1767(292)  = \1699(105)  & \1681(192) ,
  \3085(172)  = ~\3079(91) ,
  \355(399)  = \[1] ,
  \456(94)  = ~\58(7) ,
  \1971(282)  = ~\807(181) ,
  \2831(1664)  = ~\3481(1655)  | ~\3478(1653) ,
  \1025(244)  = \1022(206)  & \116(13) ,
  \3163(1181)  = \2338(1153) ,
  \1469(754)  = \1461(670)  & \322(43) ,
  \360(794)  = ~\1029(588) ,
  \2597(1509)  = ~\3393(1497)  | ~\3390(1397) ,
  \1310(597)  = ~\1099(504) ,
  \2199(1001)  = \2193(923)  & (\2173(845)  & \179(23) ),
  \989(323)  = \759(198)  & \741(116) ,
  \1027(393)  = \1024(328)  & \845(74) ,
  \1901(336)  = ~\1834(215) ,
  \2023(476)  = \807(181)  & (\274(37)  & \1817(459) ),
  \1340(808)  = \1332(646)  & \150(20) ,
  \1371(876)  = \1363(696)  & \483(81) ,
  \2077(487)  = \2076(279)  & (\250(33)  & \1799(461) ),
  \3020(163)  = \479(82) ,
  \378(1597)  = \2709(1587) ,
  \2234(480)  = \2233(278)  & (\270(36)  & \1799(461) ),
  \1742(364)  = \1739(288)  & \238(31) ,
  \1360(680)  = ~\1087(514) ,
  \1617(1356)  = ~\1616(733)  & (~\1614(1325)  & ~\1612(1127) ),
  \1283(892)  = \1275(675)  & \447(95) ,
  \1597(308)  = ~\1512(193) ,
  \1902(451)  = \1773(345)  & \1834(215) ,
  \2891(1669)  = ~\2896(1648)  | ~\2895(1659) ,
  \2143(1116)  = \2137(925)  & (\2120(1069)  & \169(22) ),
  \3277(1345)  = ~\2532(1303)  | (~\2531(1312)  | ~\2530(1141) ),
  \3491(1539)  = \2745(1521) ,
  \804(303)  = ~\776(107)  | ~\860(208) ,
  \540(65)  = ~\116(13) ,
  \1490(765)  = \1482(703)  & \303(40) ,
  \2871(128)  = \2868(50)  | \2865(61) ,
  \794(182)  = \791(103) ,
  \1612(1127)  = \1609(577)  & \1539(1079) ,
  \1458(767)  = \1450(637)  & \303(40) ,
  \1252(824)  = \1244(689)  & \137(18) ,
  \1244(689)  = ~\1123(516) ,
  \3194(1048)  = ~\3190(983) ,
  \554(219)  = \552(132)  & (\551(134)  & (\550(136)  & \549(139) )),
  \3007(97)  = \50(6) ,
  \3326(1279)  = \2433(1251) ,
  \[10]  = \383(1541)  & \2745(1521) ,
  \1636(580)  = ~\1545(470) ,
  \2978(492)  = \562(363) ,
  \2622(1422)  = ~\3418(1331)  | ~\3411(1403) ,
  \3212(1163)  = ~\3208(1139) ,
  \1379(617)  = ~\1195(507) ,
  \[11]  = \366(1577)  & \365(1570) ,
  \1066(312)  = \1057(197)  & \1049(114) ,
  \2037(1003)  = \2031(932)  & (\2013(871)  & \179(23) ),
  \2225(835)  = \2222(520)  | (\2219(380)  | \2216(740) ),
  \1087(514)  = \1084(375) ,
  \1304(810)  = \1296(708)  & \150(20) ,
  \1398(714)  = ~\1213(519) ,
  \[12]  = \386(1602)  & \2763(1589) ,
  \1604(1088)  = \1603(1031)  | \1602(1030) ,
  \1620(565)  = \1572(334)  & \1545(470) ,
  \1751(299)  = ~\1681(192) ,
  \[13]  = \392(1594)  & \2797(1582) ,
  \643(413)  = ~\3086(263)  | ~\3079(91) ,
  \393(1605)  = \[13] ,
  \1334(864)  = \1326(678)  & \492(80) ,
  \3346(1453)  = ~\3342(1427) ,
  \3419(51)  = \330(46) ,
  \3078(1121)  = ~\3074(1067) ,
  \[14]  = \389(1592)  & \2780(1580) ,
  \3193(1212)  = ~\3187(1176) ,
  \3150(1144)  = \2328(1101) ,
  \2129(484)  = \2128(276)  & (\257(34)  & \1799(461) ),
  \2204(961)  = ~\2177(846) ,
  \933(1419)  = \927(347)  & \932(1371) ,
  \1607(1033)  = \1512(193)  & \1511(911) ,
  \1474(766)  = \1466(718)  & \303(40) ,
  \1941(1123)  = ~\1916(1077) ,
  \1674(554)  = \1563(329)  & \1554(471) ,
  \714(124)  = ~\1(0) ,
  \2345(1194)  = ~\3162(1044)  | ~\3155(1180) ,
  \681(1081)  = ~\680(420)  & ~\679(1015) ,
  \1319(894)  = \1311(613)  & \447(95) ,
  \1434(652)  = ~\1231(511) ,
  \3023(268)  = ~\3017(169) ,
  \[17]  = \380(1615)  & \2728(1599) ,
  \2065(534)  = \2058(454)  & (\2052(213)  & \87(10) ),
  \3034(255)  = ~\3030(161) ,
  \[18]  = ~\406(1643) ,
  \3385(1496)  = ~\3379(1478) ,
  \2476(924)  = ~\2185(786) ,
  \399(1428)  = \[7] ,
  \[19]  = ~\408(1660) ,
  \661(1080)  = \660(274)  & \568(972) ,
  \619(1091)  = ~\2997(1038)  | ~\2994(970) ,
  \3563(1702)  = ~\3557(1695) ,
  \2577(1474)  = ~\3370(1399)  | ~\3363(1458) ,
  \3025(406)  = ~\3023(268)  | ~\3020(163) ,
  \1028(521)  = \1027(393)  | (\1026(354)  | \1025(244) ),
  \2562(1410)  = ~\3293(1379)  | ~\3290(1315) ,
  \3510(1625)  = \2690(1611) ,
  \1633(1257)  = ~\2350(1195)  | ~\2349(1232) ,
  \3478(1653)  = \2828(1640) ,
  \2409(1285)  = \2346(1256) ,
  \2354(946)  = \2013(871)  & \2289(239) ,
  \1368(847)  = \1360(680)  & \517(70) ,
  \1957(407)  = ~\1773(345)  & ~\68(8) ,
  \1259(594)  = ~\1099(504) ,
  \1987(1004)  = \1981(934)  & (\1963(881)  & \179(23) ),
  \3434(1552)  = ~\3430(1537) ,
  \2439(1281)  = \2396(1253) ,
  \1975(790)  = \1974(743)  | (\1973(477)  | \1972(493) ),
  \2888(1668)  = ~\2887(1647)  | ~\2886(1658) ,
  \3010(173)  = \456(94) ,
  \2769(560)  = ~\870(443) ,
  \2251(1000)  = \2245(920)  & (\2225(835)  & \179(23) ),
  \1632(1326)  = \1628(448)  & \1631(1286) ,
  \2848(1663)  = ~\2853(1652)  | ~\2852(1639) ,
  \665(433)  = ~\804(303) ,
  \1626(1417)  = ~\1625(732)  & (~\1623(1387)  & ~\1621(1128) ),
  \1378(601)  = ~\1186(505) ,
  \1484(639)  = ~\1222(509) ,
  \2600(1542)  = ~\2599(1527) ,
  \1023(320)  = ~\759(198) ,
  \3402(1361)  = ~\3398(1332) ,
  \2570(1491)  = ~\3361(1476)  | ~\3358(1363) ,
  \978(379)  = \975(321)  & \150(20) ,
  \[20]  = \404(1714)  & \403(1713) ,
  \2632(1415)  = ~\2629(1385) ,
  \851(68)  = ~\107(12) ,
  \1096(370)  = ~\1069(311)  | ~\1038(148) ,
  \[21]  = ~\401(1716)  | ~\400(1715) ,
  \836(85)  = ~\68(8) ,
  \3331(1516)  = \2541(1498) ,
  \3203(1213)  = ~\3197(1177) ,
  \1545(470)  = \1542(348) ,
  \1998(1112)  = \1997(1075)  & \1996(1062) ,
  \2331(1294)  = ~\3145(1268)  | ~\3142(1143) ,
  \2916(1712)  = ~\3571(1704)  | ~\3568(1694) ,
  \364(1484)  = \[8] ,
  \1799(461)  = ~\1791(344) ,
  \3525(1686)  = \2833(1681) ,
  \397(1394)  = \2657(1368)  & (\2514(1309)  & \330(46) ),
  \349(1224)  = ~\605(1186) ,
  \2395(1191)  = ~\3244(1042)  | ~\3237(1171) ,
  \3426(1344)  = ~\3422(1311) ,
  \2736(1502)  = \2733(465)  & \2581(1472) ,
  \2419(1288)  = \2359(1258) ,
  \2645(1305)  = \2467(1275) ,
  \1358(951)  = ~\1357(800)  & (~\1356(906)  & (~\1355(896)  & (~\1354(886)  & (~\1353(875)  & (~\1352(865)  & (~\1351(855)  & ~\1350(807) )))))),
  \3036(400)  = ~\3034(255)  | ~\3027(162) ,
  \1731(185)  = ~\1699(105) ,
  \3090(166)  = \898(84) ,
  \1186(505)  = \1096(370) ,
  \1584(1083)  = \1583(1021)  | \1582(1020) ,
  \3565(1696)  = \2910(1689) ,
  \2774(1572)  = \2769(560)  & \2673(1557) ,
  \1303(803)  = \1295(692)  & \159(21) ,
  \2700(1520)  = \2697(463)  & \2558(1493) ,
  \2942(57)  = \244(32) ,
  \1392(918)  = ~\1391(838)  & (~\1390(848)  & (~\1389(857)  & (~\1388(867)  & (~\1387(877)  & (~\1386(888)  & (~\1385(898)  & ~\1384(784) )))))),
  \447(95)  = \58(7) ,
  \2804(575)  = \870(443)  & \956(346) ,
  \1718(285)  = \1699(105)  & \1681(192) ,
  \398(1366)  = \2654(1337)  & \2519(1300) ,
  \1765(301)  = ~\1681(192) ,
  \635(164)  = ~\476(83)  | ~\460(89) ,
  \2677(1514)  = ~\3458(1455)  | ~\3451(1487) ,
  \1442(768)  = \1434(652)  & \303(40) ,
  \566(797)  = ~\2974(589)  | ~\2967(497) ,
  \2117(531)  = \2110(455)  & (\2052(213)  & \97(11) ),
  \1721(368)  = \1718(285)  & \223(28) ,
  \1502(656)  = ~\1231(511) ,
  \3055(532)  = ~\3036(400)  | ~\3035(394) ,
  \1663(583)  = ~\1554(471) ,
  \3490(1667)  = ~\3486(1654) ,
  \2974(589)  = ~\2970(491) ,
  \2909(1684)  = \2900(350)  & (\2892(1678)  & \2849(1673) ),
  \1318(884)  = \1310(597)  & \467(87) ,
  \1290(955)  = ~\1289(826)  & (~\1288(822)  & (~\1287(817)  & (~\1286(811)  & (~\1285(804)  & (~\1284(902)  & (~\1283(892)  & ~\1282(829) )))))),
  \941(333)  = ~\864(210) ,
  \1447(621)  = ~\1195(507) ,
  \1757(490)  = \1756(360)  | (\1755(225)  | \1754(353) ),
  \596(854)  = ~\3062(721)  | ~\3055(532) ,
  \1278(691)  = ~\1123(516) ,
  \2563(1378)  = ~\3294(1347)  | ~\3287(1346) ,
  \2332(1264)  = ~\3146(1167)  | ~\3139(1241) ,
  \3158(979)  = \2341(945) ,
  \351(1247)  = \[4] ,
  \1536(1016)  = \1533(421)  & \1256(957) ,
  \1720(235)  = \1717(183)  & \222(27) ,
  \2794(1392)  = \2787(574)  & \1671(1358) ,
  \1510(750)  = \1502(656)  & \326(44) ,
  \2586(1459)  = ~\2585(1411)  | ~\2584(1437) ,
  \1446(605)  = ~\1186(505) ,
  \3213(1240)  = \2372(1203) ,
  \1981(934)  = ~\1975(790) ,
  \2823(1631)  = ~\2822(1619)  | ~\2821(1607) ,
  \2554(1560)  = ~\2553(1531)  | ~\2552(1546) ,
  \1872(479)  = \807(181)  & (\274(37)  & \1817(459) ),
  \1393(666)  = ~\1168(513) ,
  \1388(867)  = \1380(697)  & \492(80) ,
  \1581(304)  = ~\1512(193) ,
  \657(177)  = \802(100) ,
  \552(132)  = ~\530(66)  | ~\270(36) ,
  \547(143)  = ~\467(87)  | ~\238(31) ,
  \1063(242)  = \1054(196)  & \1048(62) ,
  \2185(786)  = \2184(747)  | (\2183(473)  | \2182(483) ),
  \741(116)  = ~\20(2) ,
  \1054(196)  = \1051(112) ,
  \1862(899)  = \1859(547)  | (\1856(417)  | \1853(735) ),
  \3120(1513)  = ~\3116(1494) ,
  \2602(1449)  = ~\3402(1361)  | ~\3395(1429) ,
  \1460(914)  = ~\1459(762)  & (~\1458(767)  & (~\1457(773)  & (~\1456(780)  & (~\1455(842)  & (~\1454(852)  & (~\1453(861)  & ~\1452(758) )))))),
  \1466(718)  = ~\1213(519) ,
  \3037(157)  = \526(69) ,
  \3316(1341)  = \2426(1307) ,
  \3026(410)  = ~\3024(261)  | ~\3017(169) ,
  \2359(1258)  = ~\2358(1196)  | ~\2357(1233) ,
  \887(444)  = \867(332) ,
  \2754(1556)  = \2751(466)  & \2594(1526) ,
  \2072(863)  = ~\2065(534)  & (~\2062(395)  & ~\2059(738) ),
  \2248(1006)  = \2242(919)  & (\2225(835)  & \169(22) ),
  \479(82)  = ~\77(9) ,
  \979(543)  = \978(379)  | (\977(414)  | \976(266) ),
  \1357(800)  = \1349(647)  & \159(21) ,
  \2333(1317)  = ~\2332(1264)  | ~\2331(1294) ,
  \605(1186)  = ~\604(1159)  | ~\603(1120) ,
  \3190(983)  = \2367(947) ,
  \3174(981)  = \2354(946) ,
  \1263(626)  = ~\1147(508) ,
  \1327(598)  = ~\1099(504) ,
  \1769(221)  = \1766(190)  & \257(34) ,
  \3275(1461)  = ~\3269(1439) ,
  \861(209)  = ~\736(118)  | (~\724(119)  | ~\707(127) ),
  \2533(1193)  = ~\2454(1165) ,
  \2155(1150)  = ~\2146(1108)  & ~\2143(1116) ,
  \2379(1250)  = ~\3220(1164)  | ~\3213(1240) ,
  \1050(113)  = ~\200(25)  | ~\20(2) ,
  \2547(1545)  = ~\3337(1534)  | ~\3334(1426) ,
  \2237(785)  = \2236(748)  | (\2235(472)  | \2234(480) ),
  \2765(1590)  = ~\2760(1391)  & (~\2757(1579)  & ~\2754(1556) ),
  \1586(1022)  = \1585(305)  & \1290(955) ,
  \358(1161)  = \[3] ,
  \1730(296)  = ~\1681(192) ,
  \2868(50)  = \343(47) ,
  \2860(1710)  = ~\3540(1706)  | ~\3533(1687) ,
  \1346(695)  = ~\1123(516) ,
  \3403(1402)  = \2609(1369) ,
  \1947(1170)  = \1946(1146)  & \1945(1155) ,
  \950(1547)  = ~\955(1536)  | ~\954(1532) ,
  \1661(1126)  = \1656(552)  & \673(1082) ,
  \2751(466)  = ~\956(346) ,
  \1269(818)  = \1261(690)  & \143(19) ,
  \2042(964)  = ~\2017(872) ,
  \3259(1383)  = ~\3253(1352) ,
  \736(118)  = \20(2) ,
  \1465(702)  = ~\1204(517) ,
  \1377(681)  = ~\1177(515) ,
  \2678(462)  = ~\956(346) ,
  \560(226)  = ~\2945(142)  | ~\2942(57) ,
  \1002(317)  = ~\759(198) ,
  \590(891)  = ~\3054(726)  | ~\3047(546) ,
  \3070(1119)  = ~\3066(1066) ,
  \396(1504)  = \[9] ,
  \1939(1105)  = \1930(936)  & (\1916(1077)  & \190(24) ),
  \3179(1179)  = \2351(1152) ,
  \1123(516)  = \1120(376) ,
  \1639(1130)  = \1636(580)  & \1592(1085) ,
  \1111(506)  = \1108(371) ,
  \1613(1293)  = ~\1615(1263) ,
  \654(256)  = ~\626(158)  | ~\87(10) ,
  \3494(1627)  = \2839(1614) ,
  \3337(1534)  = ~\3331(1516) ,
  \704(126)  = ~\1(0) ,
  \3547(1645)  = ~\3541(1632) ,
  \997(259)  = \994(202)  & \77(9) ,
  \3524(1671)  = ~\3520(1661) ,
  \3438(1500)  = \2638(1483) ,
  \2102(1071)  = \2099(963)  | (\2098(989)  | \2097(995) ),
  \555(231)  = ~\2937(146)  | ~\2934(59) ,
  \2837(1675)  = ~\3490(1667)  | ~\3483(1642) ,
  \1247(641)  = ~\1159(510) ,
  \2917(1703)  = ~\3572(1700)  | ~\3565(1696) ,
  \780(106)  = ~\33(3) ,
  \2285(241)  = \213(26)  & \2278(207) ,
  \2209(1068)  = \2204(961)  | (\2203(988)  | \2202(994) ),
  \1007(528)  = \1006(409)  | (\1005(392)  | \1004(252) ),
  \3532(1705)  = ~\3528(1697) ,
  \1621(1128)  = \1618(578)  & \1584(1083) ,
  \2680(568)  = \870(443)  & \956(346) ,
  \992(418)  = \989(323)  & \50(6) ,
  \1177(515)  = \1084(375) ,
  \2386(1227)  = ~\3235(1211)  | ~\3232(976) ,
  \1461(670)  = ~\1168(513) ,
  \1991(991)  = \1978(933)  & (\1967(882)  & \200(25) ),
  \3319(1367)  = ~\3313(1336) ,
  \1960(540)  = \1953(452)  & (\1829(214)  & \68(8) ),
  \562(363)  = ~\561(229)  | ~\560(226) ,
  \1681(192)  = \780(106) ,
  \1601(309)  = ~\1512(193) ,
  \3355(1457)  = \2564(1435) ,
  \2505(1320)  = \2268(1245)  & \2495(1283) ,
  \1794(460)  = \1791(344) ,
  \1893(1064)  = ~\1886(1005)  & ~\1883(1011) ,
  \3430(1537)  = \2635(1465)  & \2572(1510) ,
  \557(366)  = ~\556(233)  | ~\555(231) ,
  \3216(1140)  = \2375(1097) ,
  \1338(905)  = \1330(710)  & \432(99) ,
  \1402(889)  = \1394(682)  & \467(87) ,
  \3329(1162)  = ~\3323(1138) ,
  \3572(1700)  = ~\3568(1694) ,
  \641(728)  = \639(272)  & (\476(83)  & \640(541) ),
  \1445(685)  = ~\1177(515) ,
  \1606(1032)  = \1605(310)  & \1375(950) ,
  \3474(1618)  = ~\3470(1601) ,
  \2183(473)  = \816(179)  & (\274(37)  & \1799(461) ),
  \3229(1174)  = \2380(1148) ,
  \842(77)  = ~\87(10) ,
  \2378(1278)  = ~\3219(1267)  | ~\3216(1140) ,
  \2308(1271)  = ~\2275(1246) ,
  \2028(931)  = \2025(789) ,
  \405(1717)  = \[20] ,
  \354(257)  = \626(158)  & \87(10) ,
  \995(316)  = ~\759(198) ,
  \1642(1259)  = ~\2363(1197)  | ~\2362(1234) ,
  \1459(762)  = \1451(653)  & \311(41) ,
  \1373(897)  = \1365(632)  & \447(95) ,
  \2663(1567)  = \2662(1548)  | \2661(1561) ,
  \1331(630)  = ~\1147(508) ,
  \2986(355)  = ~\2966(220)  | ~\2965(218) ,
  \1132(377)  = ~\1060(243)  | ~\1043(149) ,
  \625(167)  = \836(85)  & (\831(92)  & \826(96) ),
  \1637(449)  = ~\1572(334) ,
  \913(390)  = ~\3110(251)  | ~\3103(71) ,
  \2816(1468)  = ~\2811(1393)  & (~\2808(1443)  & ~\2805(1446) ),
  \2556(1475)  = ~\3353(1456)  | ~\3350(1334) ,
  \1505(770)  = \1497(608)  & \294(39) ,
  \1641(1327)  = \1637(449)  & \1640(1289) ,
  \2013(871)  = \2010(537)  | (\2007(401)  | \2004(737) ),
  \3050(539)  = ~\3026(410)  | ~\3025(406) ,
  \3145(1268)  = ~\3139(1241) ,
  \1475(761)  = \1467(638)  & \311(41) ,
  \1748(228)  = \1745(187)  & \238(31) ,
  \634(247)  = ~\905(155)  | ~\540(65) ,
  \1351(855)  = \1343(679)  & \504(76) ,
  \1722(502)  = \1721(368)  | (\1720(235)  | \1719(402) ),
  \1222(509)  = \1144(372) ,
  \1315(645)  = ~\1159(510) ,
  \579(939)  = \576(793) ,
  \1770(357)  = \1767(292)  & \264(35) ,
  \2703(1578)  = \2698(556)  & \2666(1565) ,
  \1308(661)  = ~\1075(512) ,
  \1923(742)  = \1729(501)  & \1812(458) ,
  \1414(699)  = ~\1204(517) ,
  \2908(1676)  = \2903(349)  & (\2888(1668)  & \2849(1673) ),
  \3024(261)  = ~\3020(163) ,
  \3370(1399)  = ~\3366(1364) ,
  \1390(848)  = \1382(633)  & \517(70) ,
  \1610(446)  = ~\1572(334) ,
  \1486(751)  = \1478(671)  & \326(44) ,
  \2080(788)  = \2079(745)  | (\2078(475)  | \2077(487) ),
  \3409(1430)  = ~\3403(1402) ,
  \2900(350)  = \2897(49)  & \2877(217) ,
  \1011(909)  = \1008(204)  & \911(724) ,
  \1240(657)  = ~\1075(512) ,
  \1759(189)  = ~\1699(105) ,
  \1491(760)  = \1483(719)  & \311(41) ,
  \2003(453)  = \1773(345)  & \1834(215) ,
  \976(266)  = \973(199)  & \897(168) ,
  \3390(1397)  = \2589(1362) ,
  \1754(353)  = \1751(299)  & \283(38) ,
  \2929(1644)  = \2925(1629)  & \2922(1608) ,
  \1664(438)  = ~\1563(329) ,
  \3564(1699)  = ~\3560(1693) ,
  \671(426)  = ~\806(293) ,
  \604(1159)  = ~\3078(1121)  | ~\3071(1014) ,
  \2078(475)  = \823(180)  & (\274(37)  & \1799(461) ),
  \1396(618)  = ~\1195(507) ,
  \2684(1596)  = \2679(555)  & \2660(1584) ,
  \3462(1593)  = \2797(1582) ,
  \2235(472)  = \816(179)  & (\274(37)  & \1799(461) ),
  \1634(730)  = \1629(566)  & \463(88) ,
  \2763(1589)  = \2760(1391)  | (\2757(1579)  | \2754(1556) ),
  \2998(1036)  = ~\2994(970) ,
  \2609(1369)  = ~\2608(1339)  | ~\2607(1301) ,
  \2821(1607)  = ~\3465(1505)  | ~\3462(1593) ,
  \2673(1557)  = ~\2672(1524)  | ~\2671(1550) ,
  \2945(142)  = ~\2939(58) ,
  \2808(1443)  = \2803(562)  & \2626(1395) ,
  \2535(1338)  = ~\2461(1137)  | (~\2433(1251)  | ~\2426(1307) ),
  \731(121)  = \20(2)  & \13(1) ,
  \2989(486)  = ~\2983(359) ,
  \915(331)  = ~\861(209) ,
  \381(1626)  = \[17] ,
  \1984(1010)  = \1978(933)  & (\1963(881)  & \169(22) ),
  \2753(572)  = \870(443)  & \956(346) ,
  \2152(1149)  = \2146(1108)  | \2143(1116) ,
  \662(550)  = \657(177)  & \655(416) ,
  \1477(913)  = ~\1476(757)  & (~\1475(761)  & (~\1474(766)  & (~\1473(772)  & (~\1472(779)  & (~\1471(843)  & (~\1470(853)  & ~\1469(754) )))))),
  \636(175)  = \442(98) ,
  \1253(828)  = \1245(705)  & \132(17) ,
  \3248(978)  = \2391(944) ,
  \2425(1249)  = ~\3212(1163)  | ~\3205(1239) ,
  \791(103)  = ~\41(4) ,
  \3171(1178)  = \2351(1152) ,
  \1372(887)  = \1364(712)  & \467(87) ,
  \2852(1639)  = ~\3505(1555)  | ~\3502(1628) ,
  \1669(1252)  = ~\2387(1190)  | ~\2386(1227) ,
  \1451(653)  = ~\1231(511) ,
  \1305(816)  = \1297(628)  & \143(19) ,
  \2477(921)  = ~\2237(785) ,
  \2002(338)  = ~\1834(215) ,
  \2635(1465)  = ~\2634(1416)  & ~\2633(1420) ,
  \655(416)  = \58(7)  & (\442(98)  & (\635(164)  & \630(246) )),
  \3450(1515)  = ~\3446(1495) ,
  \1668(1323)  = \1664(438)  & \1667(1280) ,
  \2315(1244)  = ~\2314(1205)  | (~\2313(1209)  | (~\2312(1175)  | ~\2311(1109) )),
  \890(125)  = \1(0) ,
  \526(69)  = ~\107(12) ,
  \2193(923)  = ~\2185(786) ,
  \363(1466)  = ~\1030(1442) ,
  \1031(1571)  = ~\951(1564)  & (~\947(910)  & ~\944(969) ),
  \3295(1276)  = \2464(1248) ,
  \1660(1308)  = ~\2379(1250)  | ~\2378(1278) ,
  \1276(595)  = ~\1099(504) ,
  \1395(602)  = ~\1186(505) ,
  \3243(1207)  = ~\3237(1171) ,
  \3014(271)  = ~\3010(173) ,
  \1595(1027)  = \1512(193)  & \1460(914) ,
  \2713(1588)  = ~\2706(1444)  & (~\2703(1578)  & ~\2700(1520) ),
  \2458(1096)  = \2302(236)  & \2257(1053) ,
  \1967(882)  = ~\1960(540)  & (~\1957(407)  & ~\1954(736) ),
  \3074(1067)  = \600(1012) ,
  \3483(1642)  = \2823(1631) ,
  \1335(874)  = \1327(598)  & \483(81) ,
  \2101(1058)  = ~\2094(1002)  & ~\2091(1008) ,
  \2786(561)  = ~\870(443) ,
  \1389(857)  = \1381(713)  & \504(76) ,
  \2254(993)  = \2245(920)  & (\2229(836)  & \190(24) ),
  \3342(1427)  = \2544(1400) ,
  \2842(1638)  = ~\3497(1554)  | ~\3494(1627) ,
  \2097(995)  = \2088(929)  & (\2072(863)  & \190(24) ),
  \2491(1255)  = \2490(1230)  | \2489(1100) ,
  \2768(467)  = ~\956(346) ,
  \3556(1622)  = ~\3552(1610) ,
  \2132(787)  = \2131(746)  | (\2130(474)  | \2129(484) ),
  \1024(328)  = \759(198)  & \741(116) ,
  \2576(1492)  = ~\3369(1477)  | ~\3366(1364) ,
  \2981(592)  = ~\2975(498) ,
  \3427(1512)  = \2558(1493) ,
  \2261(1065)  = \2256(959)  | (\2255(987)  | \2254(993) ),
  \620(1093)  = ~\2998(1036)  | ~\2991(973) ,
  \644(269)  = \636(175)  & \460(89) ,
  \1572(334)  = ~\784(191)  | ~\724(119) ,
  \2621(1448)  = ~\3417(1431)  | ~\3414(1298) ,
  \1419(879)  = \1411(683)  & \483(81) ,
  \3169(1220)  = ~\3163(1181) ,
  \3094(265)  = ~\3090(166) ,
  \2265(1215)  = \2048(1111)  & (\1998(1112)  & (\1947(1170)  & \1895(1115) )),
  \3131(1184)  = \2317(1156) ,
  \3121(1183)  = \2317(1156) ,
  \3221(1173)  = \2380(1148) ,
  \1375(950)  = ~\1374(907)  & (~\1373(897)  & (~\1372(887)  & (~\1371(876)  & (~\1370(866)  & (~\1369(856)  & (~\1368(847)  & ~\1367(799) )))))),
  \3016(419)  = ~\3014(271)  | ~\3007(97) ,
  \2650(1404)  = \2647(1372) ,
  \660(274)  = ~\657(177) ,
  \1248(834)  = \1240(657)  & \124(14) ,
  \1635(1355)  = ~\1634(730)  & (~\1632(1326)  & ~\1630(1129) ),
  \2589(1362)  = \2513(1343)  & \330(46) ,
  \994(202)  = ~\741(116) ,
  \3414(1298)  = \2612(1272) ,
  \2275(1246)  = ~\2274(1214)  | (~\2273(1218)  | (~\2272(1182)  | ~\2271(1114) )),
  \1015(205)  = ~\741(116) ,
  \2448(1099)  = \2293(238)  & \2043(1059) ,
  \2514(1309)  = \2433(1251)  & \2439(1281) ,
  \1540(111)  = ~\20(2) ,
  \3027(162)  = \501(79) ,
  \367(1585)  = \[11] ,
  \1295(692)  = ~\1123(516) ,
  \3269(1439)  = \2527(1412) ,
  \3320(1374)  = ~\3316(1341) ,
  \2629(1385)  = \2501(1353) ,
  \690(535)  = \685(427)  & \654(256) ,
  \1749(362)  = \1746(289)  & \244(32) ,
  \3113(1499)  = ~\3112(1464)  | ~\3111(1482) ,
  \1993(1061)  = \1987(1004)  | \1984(1010) ,
  \2928(1623)  = \2874(129)  & (\2694(1612)  & \2713(1588) ),
  \639(272)  = ~\636(175) ,
  \1464(622)  = ~\1195(507) ,
  \3252(1043)  = ~\3248(978) ,
  \3506(1637)  = ~\3502(1628) ,
  \1478(671)  = ~\1168(513) ,
  \2482(949)  = \2481(150)  & (\2237(785)  & (\2185(786)  & (\2132(787)  & \2080(788) ))),
  \548(141)  = ~\483(81)  | ~\244(32) ,
  \614(968)  = \610(432)  & \576(793) ,
  \1651(1261)  = ~\2371(1199)  | ~\2370(1236) ,
  \2088(929)  = ~\2080(788) ,
  \974(313)  = ~\759(198) ,
  \1648(1131)  = \1645(581)  & \1596(1086) ,
  \2451(1142)  = \2448(1099) ,
  \3457(1506)  = ~\3451(1487) ,
  \3232(976)  = \2383(943) ,
  \1213(519)  = \1132(377) ,
  \1316(820)  = \1308(661)  & \137(18) ,
  \2245(920)  = ~\2237(785) ,
  \1973(477)  = \807(181)  & (\274(37)  & \1817(459) ),
  \2676(1533)  = ~\3457(1506)  | ~\3454(1432) ,
  \1746(289)  = \1699(105)  & \1681(192) ,
  \1877(937)  = \1874(792) ,
  \3061(725)  = ~\3055(532) ,
  \2461(1137)  = \2458(1096) ,
  \1630(1129)  = \1627(579)  & \1588(1084) ,
  \3129(1237)  = ~\3127(1221)  | ~\3124(985) ,
  \1627(579)  = ~\1545(470) ,
  \833(86)  = \68(8) ,
  \669(1019)  = \665(433)  & \597(960) ,
  \3161(1219)  = ~\3155(1180) ,
  \3322(1401)  = ~\3320(1374)  | ~\3313(1336) ,
  \1483(719)  = ~\1213(519) ,
  \1512(193)  = \776(107) ,
  \513(75)  = ~\97(11) ,
  \1593(307)  = ~\1512(193) ,
  \2624(1329)  = ~\3425(130)  | ~\3422(1311) ,
  \1658(1342)  = ~\1660(1308) ,
  \1638(567)  = \1572(334)  & \1545(470) ,
  \1891(967)  = ~\1866(900) ,
  \3358(1363)  = \2567(1333) ,
  \3374(1273)  = \2491(1255)  & \330(46) ,
  \1348(631)  = ~\1147(508) ,
  \3063(1013)  = \591(965) ,
  \3507(1598)  = \2709(1587) ,
  \1738(186)  = ~\1699(105) ,
  \568(972)  = ~\567(941) ,
  \893(216)  = \890(125) ,
  \1892(1063)  = \1886(1005)  | \1883(1011) ,
  \2501(1353)  = \2500(1319)  | \2275(1246) ,
  \1051(112)  = \179(23)  & \20(2) ,
  \3220(1164)  = ~\3216(1140) ,
  \404(1714)  = ~\2917(1703)  | ~\2916(1712) ,
  \1286(811)  = \1278(691)  & \150(20) ,
  \1280(627)  = ~\1147(508) ,
  \2363(1197)  = ~\3186(1047)  | ~\3179(1179) ,
  \3139(1241)  = \2325(1204) ,
  \2865(61)  = ~\213(26) ,
  \2481(150)  = ~\2478(64) ,
  \1344(599)  = ~\1099(504) ,
  \2822(1619)  = ~\3466(1606)  | ~\3459(1485) ,
  \3162(1044)  = ~\3158(979) ,
  \2151(1122)  = ~\2124(1070) ,
  \2271(1114)  = ~\1892(1063) ,
  \2307(1270)  = ~\2315(1244)  | ~\2265(1215) ,
  \350(1223)  = ~\608(1185) ,
  \1463(606)  = ~\1186(505) ,
  \679(1015)  = \678(275)  & \591(965) ,
  \2922(1608)  = \2765(1590)  & (\2782(1581)  & (\2799(1583)  & \2816(1468) )),
  \3571(1704)  = ~\3565(1696) ,
  \3486(1654)  = \2828(1640) ,
  \2489(1100)  = \2488(503)  & \2484(1052) ,
  \2262(1106)  = \2261(1065)  & \2260(1054) ,
  \1394(682)  = ~\1177(515) ,
  \3393(1497)  = ~\3387(1479) ,
  \3106(154)  = \907(67) ,
  \561(229)  = ~\2946(140)  | ~\2939(58) ,
  \2047(1072)  = \2042(964)  | (\2041(990)  | \2040(996) ),
  \2130(474)  = \816(179)  & (\274(37)  & \1799(461) ),
  \1403(878)  = \1395(602)  & \483(81) ,
  \1650(1322)  = \1646(436)  & \1649(1291) ,
  \2364(1151)  = \2103(1110) ,
  \1766(190)  = ~\1699(105) ,
  \1482(703)  = ~\1204(517) ,
  \2068(862)  = \2065(534)  | (\2062(395)  | \2059(738) ),
  \973(199)  = ~\741(116) ,
  \1852(450)  = \1773(345)  & \1834(215) ,
  \3523(1680)  = ~\3517(1672) ,
  \1936(1113)  = \1930(936)  & (\1912(1076)  & \179(23) ),
  \476(83)  = \77(9) ,
  \1945(1155)  = ~\1936(1113)  & ~\1933(1117) ,
  \923(482)  = \916(442)  & \586(356) ,
  \1257(658)  = ~\1075(512) ,
  \2208(1056)  = ~\2199(1001)  & ~\2196(1007) ,
  \2910(1689)  = \2909(1684)  | (\2908(1676)  | (\2907(1683)  | \2906(1677) )),
  \606(1118)  = ~\3069(1073)  | ~\3066(1066) ,
  \2444(1166)  = \2288(240)  & \1942(1154) ,
  \2454(1165)  = \2293(238)  & \2152(1149) ,
  \688(428)  = \806(293)  & \804(303) ,
  \2839(1614)  = \2728(1599) ,
  \1003(325)  = \759(198)  & \741(116) ,
  \947(910)  = \942(441)  & \649(723) ,
  \517(70)  = \107(12) ,
  \2534(1335)  = ~\2455(1095)  | ~\2426(1307) ,
  \977(414)  = \974(313)  & \828(93) ,
  \996(324)  = \759(198)  & \741(116) ,
  \1264(642)  = ~\1159(510) ,
  \556(233)  = ~\2938(144)  | ~\2931(60) ,
  \1592(1085)  = \1591(1025)  | \1590(1024) ,
  \1649(1291)  = ~\1651(1261) ,
  \2464(1248)  = \2302(236)  & \2315(1244) ,
  \2864(1709)  = ~\3532(1705)  | ~\3525(1686) ,
  \2024(744)  = \1743(496)  & \1812(458) ,
  \1416(635)  = ~\1222(509) ,
  \3533(1687)  = \2833(1681) ,
  \2344(1231)  = ~\3161(1219)  | ~\3158(979) ,
  \2388(1147)  = \2262(1106) ,
  \1728(367)  = \1725(286)  & \226(29) ,
  \1727(234)  = \1724(184)  & \223(28) ,
  \806(293)  = ~\780(106)  | ~\860(208) ,
  \1468(654)  = ~\1231(511) ,
  \1506(764)  = \1498(624)  & \303(40) ,
  \1851(335)  = ~\1834(215) ,
  \366(1577)  = ~\1031(1571) ,
  \1285(804)  = \1277(611)  & \159(21) ,
  \1906(411)  = ~\1773(345)  & ~\58(7) ,
  \1665(553)  = \1563(329)  & \1554(471) ,
  \3200(984)  = \2367(947) ,
  \1363(696)  = ~\1123(516) ,
  \380(1615)  = ~\2730(1600) ,
  \2527(1412)  = ~\2526(1370)  | (~\2525(1377)  | (~\2524(1375)  | ~\2523(1200) )),
  \1611(564)  = \1572(334)  & \1545(470) ,
  \1391(838)  = \1383(649)  & \530(66) ,
  \2836(1666)  = ~\3489(1656)  | ~\3486(1654) ,
  \1631(1286)  = ~\1633(1257) ;
endmodule

