// IWLS benchmark module "C2670.iscas" printed on Wed May 29 16:27:57 2002
module test2 (\1(0) , \2(1) , \3(2) , \4(3) , \5(4) , \6(5) , \7(6) , \8(7) ,
 \11(8) , \14(9) , \15(10) , \16(11) , \19(12) , \20(13) , \21(14) , \22(15) ,
 \23(16) , \24(17) , \25(18) , \26(19) , \27(20) , \28(21) , \29(22) , \32(23) ,
 \33(24) , \34(25) , \35(26) , \36(27) , \37(28) , \40(29) , \43(30) , \44(31) ,
 \47(32) , \48(33) , \49(34) , \50(35) , \51(36) , \52(37) , \53(38) , \54(39) ,
 \55(40) , \56(41) , \57(42) , \60(43) , \61(44) , \62(45) , \63(46) , \64(47) ,
 \65(48) , \66(49) , \67(50) , \68(51) , \69(52) , \72(53) , \73(54) , 
\74(55) , \75(56) , \76(57) , \77(58) , \78(59) , \79(60) , \80(61) , 
\81(62) , \82(63) , \85(64) , \86(65) , \87(66) , \88(67) , \89(68) , 
\90(69) , \91(70) , \92(71) , \93(72) , \94(73) , \95(74) , \96(75) , 
\99(76) , \100(77) , \101(78) , \102(79) , \103(80) , \104(81) , 
\105(82) , \106(83) , \107(84) , \108(85) , \111(86) , \112(87) , 
\113(88) , \114(89) , \115(90) , \116(91) , \117(92) , \118(93) , 
\119(94) , \120(95) , \123(96) , \124(97) , \125(98) , \126(99) , 
\127(100) , \128(101) , \129(102) , \130(103) , \131(104) , \132(105) , 
\135(106) , \136(107) , \137(108) , \138(109) , \139(110) , \140(111) , 
\141(112) , \142(113) , \IN-169(114) , \IN-174(115) , \IN-177(116) , 
\IN-178(117) , \IN-179(118) , \IN-180(119) , \IN-181(120) , \IN-182(121) , 
\IN-183(122) , \IN-184(123) , \IN-185(124) , \IN-186(125) , \IN-189(126) , 
\IN-190(127) , \IN-191(128) , \IN-192(129) , \IN-193(130) , \IN-194(131) , 
\IN-195(132) , \IN-196(133) , \IN-197(134) , \IN-198(135) , \IN-199(136) , 
\IN-200(137) , \IN-201(138) , \IN-202(139) , \IN-203(140) , \IN-204(141) , 
\IN-205(142) , \IN-206(143) , \IN-207(144) , \IN-208(145) , \IN-209(146) , 
\IN-210(147) , \IN-211(148) , \IN-212(149) , \IN-213(150) , \IN-214(151) , 
\IN-215(152) , \IN-239(153) , \IN-240(154) , \IN-241(155) , \IN-242(156) , 
\IN-243(157) , \IN-244(158) , \IN-245(159) , \IN-246(160) , \IN-247(161) , 
\IN-248(162) , \IN-249(163) , \IN-250(164) , \IN-251(165) , \IN-252(166) , 
\IN-253(167) , \IN-254(168) , \IN-255(169) , \IN-256(170) , \IN-257(171) , 
\IN-262(172) , \IN-263(173) , \IN-264(174) , \IN-265(175) , \IN-266(176) , 
\IN-267(177) , \IN-268(178) , \IN-269(179) , \IN-270(180) , \IN-271(181) , 
\IN-272(182) , \IN-273(183) , \IN-274(184) , \IN-275(185) , \IN-276(186) , 
\IN-277(187) , \IN-278(188) , \IN-279(189) , \452(190) , \483(191) , 
\543(192) , \559(193) , \567(194) , \651(195) , \661(196) , \860(197) , 
\868(198) , \1083(199) , \1341(200) , \1348(201) , \1384(202) , \1956(203) , 
\1961(204) , \1966(205) , \1971(206) , \1976(207) , \1981(208) , \1986(209) , 
\1991(210) , \1996(211) , \2066(212) , \2067(213) , \2072(214) , \2078(215) , 
\2084(216) , \2090(217) , \2096(218) , \2100(219) , \2104(220) , \2105(221) , 
\2106(222) , \2427(223) , \2430(224) , \2435(225) , \2438(226) , \2443(227) , 
\2446(228) , \2451(229) , \2454(230) , \2474(231) , \2678(232) , \169(114) , 
\174(115) , \177(116) , \178(117) , \179(118) , \180(119) , \181(120) , 
\182(121) , \183(122) , \184(123) , \185(124) , \186(125) , \189(126) , 
\190(127) , \191(128) , \192(129) , \193(130) , \194(131) , \195(132) , 
\196(133) , \197(134) , \198(135) , \199(136) , \200(137) , \201(138) , 
\202(139) , \203(140) , \204(141) , \205(142) , \206(143) , \207(144) , 
\208(145) , \209(146) , \210(147) , \211(148) , \212(149) , \213(150) , 
\214(151) , \215(152) , \239(153) , \240(154) , \241(155) , \242(156) , 
\243(157) , \244(158) , \245(159) , \246(160) , \247(161) , \248(162) , 
\249(163) , \250(164) , \251(165) , \252(166) , \253(167) , \254(168) , 
\255(169) , \256(170) , \257(171) , \262(172) , \263(173) , \264(174) , 
\265(175) , \266(176) , \267(177) , \268(178) , \269(179) , \270(180) , 
\271(181) , \272(182) , \273(183) , \274(184) , \275(185) , \276(186) , 
\277(187) , \278(188) , \279(189) , \350(301) , \335(299) , \409(298) , 
\369(289) , \367(288) , \411(264) , \337(263) , \384(262) , \218(311) , 
\219(302) , \220(306) , \221(305) , \235(307) , \236(303) , \237(309) , 
\238(304) , \158(349) , \259(414) , \391(379) , \173(389) , \223(413) , 
\234(376) , \217(423) , \325(507) , \261(506) , \319(656) , \160(609) , 
\162(612) , \164(607) , \166(625) , \168(623) , \171(621) , \153(671) , 
\176(803) , \188(761) , \299(692) , \301(694) , \286(696) , \303(698) , 
\288(700) , \305(702) , \290(704) , \284(847) , \321(848) , \297(849) , 
\280(850) , \148(851) , \282(922) , \323(923) , \156(1046) , \401(1276) , 
\227(1179) , \229(1180) , \311(1278) , \150(1277) , \145(1358) , 
\395(1392) , \295(1400) , \331(1401) , \397(1406) , \329(1414) , 
\231(1422) , \308(1425) , \225(1424) );
input
  \124(97) ,
  \IN-177(116) ,
  \111(86) ,
  \IN-239(153) ,
  \IN-174(115) ,
  \69(52) ,
  \56(41) ,
  \43(30) ,
  \IN-207(144) ,
  \1348(201) ,
  \102(79) ,
  \93(72) ,
  \IN-276(186) ,
  \14(9) ,
  \80(61) ,
  \452(190) ,
  \IN-273(183) ,
  \128(101) ,
  \2454(230) ,
  \115(90) ,
  \IN-204(141) ,
  \47(32) ,
  \34(25) ,
  \21(14) ,
  \IN-185(124) ,
  \IN-252(166) ,
  \119(94) ,
  \106(83) ,
  \IN-215(152) ,
  \25(18) ,
  \1986(209) ,
  \IN-271(181) ,
  \IN-199(136) ,
  \IN-266(176) ,
  \1083(199) ,
  \88(67) ,
  \75(56) ,
  \IN-263(173) ,
  \62(45) ,
  \IN-250(164) ,
  \IN-178(117) ,
  \29(22) ,
  \2(1) ,
  \16(11) ,
  \IN-208(145) ,
  \IN-242(156) ,
  \66(49) ,
  \53(38) ,
  \2066(212) ,
  \129(102) ,
  \79(60) ,
  \40(29) ,
  \IN-277(187) ,
  \IN-205(142) ,
  \IN-274(184) ,
  \4(3) ,
  \1981(208) ,
  \90(69) ,
  \IN-189(126) ,
  \125(98) ,
  \112(87) ,
  \IN-240(154) ,
  \1976(207) ,
  \6(5) ,
  \IN-256(170) ,
  \57(42) ,
  \44(31) ,
  \IN-253(167) ,
  \94(73) ,
  \8(7) ,
  \81(62) ,
  \116(91) ,
  \139(110) ,
  \559(193) ,
  \103(80) ,
  \IN-267(177) ,
  \48(33) ,
  \IN-251(165) ,
  \IN-264(174) ,
  \35(26) ,
  \22(15) ,
  \2072(214) ,
  \IN-179(118) ,
  \85(64) ,
  \72(53) ,
  \1971(206) ,
  \IN-246(160) ,
  \107(84) ,
  \543(192) ,
  \IN-243(157) ,
  \135(106) ,
  \2067(213) ,
  \26(19) ,
  \2435(225) ,
  \IN-209(146) ,
  \IN-278(188) ,
  \IN-275(185) ,
  \89(68) ,
  \1966(205) ,
  \76(57) ,
  \63(46) ,
  \50(35) ,
  \2078(215) ,
  \2451(229) ,
  \IN-192(129) ,
  \IN-241(155) ,
  \IN-257(171) ,
  \2446(228) ,
  \IN-254(168) ,
  \IN-169(114) ,
  \130(103) ,
  \54(39) ,
  \67(50) ,
  \11(8) ,
  \2430(224) ,
  \IN-190(127) ,
  \IN-268(178) ,
  \126(99) ,
  \2678(232) ,
  \IN-265(175) ,
  \91(70) ,
  \1961(204) ,
  \113(88) ,
  \100(77) ,
  \1956(203) ,
  \860(197) ,
  \32(23) ,
  \IN-247(161) ,
  \IN-182(121) ,
  \136(107) ,
  \IN-244(158) ,
  \95(74) ,
  \140(111) ,
  \82(63) ,
  \104(81) ,
  \IN-279(189) ,
  \IN-212(149) ,
  \IN-196(133) ,
  \49(34) ,
  \2084(216) ,
  \117(92) ,
  \36(27) ,
  \23(16) ,
  \IN-180(119) ,
  \99(76) ,
  \86(65) ,
  \73(54) ,
  \IN-193(130) ,
  \60(43) ,
  \108(85) ,
  \2104(220) ,
  \IN-255(169) ,
  \131(104) ,
  \IN-210(147) ,
  \27(20) ,
  \77(58) ,
  \1(0) ,
  \64(47) ,
  \51(36) ,
  \IN-191(128) ,
  \IN-269(179) ,
  \IN-202(139) ,
  \IN-186(125) ,
  \3(2) ,
  \IN-183(122) ,
  \IN-248(162) ,
  \661(196) ,
  \123(96) ,
  \141(112) ,
  \2090(217) ,
  \68(51) ,
  \IN-245(159) ,
  \137(108) ,
  \55(40) ,
  \5(4) ,
  \IN-200(137) ,
  \1384(202) ,
  \IN-197(134) ,
  \114(89) ,
  \2474(231) ,
  \1341(200) ,
  \92(71) ,
  \IN-213(150) ,
  \101(78) ,
  \1996(211) ,
  \7(6) ,
  \IN-181(120) ,
  \IN-194(131) ,
  \2096(218) ,
  \33(24) ,
  \20(13) ,
  \483(191) ,
  \2105(221) ,
  \567(194) ,
  \132(105) ,
  \96(75) ,
  \IN-211(148) ,
  \IN-206(143) ,
  \118(93) ,
  \105(82) ,
  \37(28) ,
  \24(17) ,
  \127(100) ,
  \IN-272(182) ,
  \87(66) ,
  \IN-203(140) ,
  \651(195) ,
  \74(55) ,
  \61(44) ,
  \1991(210) ,
  \2427(223) ,
  \IN-249(163) ,
  \IN-184(123) ,
  \142(113) ,
  \2443(227) ,
  \138(109) ,
  \28(21) ,
  \120(95) ,
  \15(10) ,
  \78(59) ,
  \IN-201(138) ,
  \65(48) ,
  \52(37) ,
  \IN-198(135) ,
  \IN-270(180) ,
  \IN-214(151) ,
  \2438(226) ,
  \2100(219) ,
  \IN-195(132) ,
  \IN-262(172) ,
  \868(198) ,
  \2106(222) ,
  \19(12) ;
output
  \269(179) ,
  \215(152) ,
  \156(1046) ,
  \397(1406) ,
  \180(119) ,
  \145(1358) ,
  \191(128) ,
  \200(137) ,
  \186(125) ,
  \197(134) ,
  \242(156) ,
  \264(174) ,
  \211(148) ,
  \206(143) ,
  \253(167) ,
  \275(185) ,
  \248(162) ,
  \311(1278) ,
  \367(288) ,
  \301(694) ,
  \225(1424) ,
  \401(1276) ,
  \181(120) ,
  \391(379) ,
  \270(180) ,
  \162(612) ,
  \192(129) ,
  \350(301) ,
  \201(138) ,
  \243(157) ,
  \265(175) ,
  \198(135) ,
  \212(149) ,
  \207(144) ,
  \254(168) ,
  \249(163) ,
  \168(623) ,
  \284(847) ,
  \150(1277) ,
  \276(186) ,
  \319(656) ,
  \261(506) ,
  \299(692) ,
  \288(700) ,
  \295(1400) ,
  \384(262) ,
  \182(121) ,
  \193(130) ,
  \271(181) ,
  \164(607) ,
  \219(302) ,
  \335(299) ,
  \235(307) ,
  \202(139) ,
  \177(116) ,
  \244(158) ,
  \239(153) ,
  \208(145) ,
  \255(169) ,
  \218(311) ,
  \199(136) ,
  \266(176) ,
  \277(187) ,
  \323(923) ,
  \369(289) ,
  \282(922) ,
  \303(698) ,
  \409(298) ,
  \183(122) ,
  \250(164) ,
  \234(376) ,
  \272(182) ,
  \194(131) ,
  \321(848) ,
  \203(140) ,
  \337(263) ,
  \256(170) ,
  \236(303) ,
  \229(1180) ,
  \259(414) ,
  \325(507) ,
  \178(117) ,
  \245(159) ,
  \176(803) ,
  \189(126) ,
  \153(671) ,
  \267(177) ,
  \329(1414) ,
  \209(146) ,
  \278(188) ,
  \213(150) ,
  \188(761) ,
  \231(1422) ,
  \220(306) ,
  \160(609) ,
  \297(849) ,
  \240(154) ,
  \184(123) ,
  \251(165) ,
  \195(132) ,
  \262(172) ,
  \273(183) ,
  \204(141) ,
  \217(423) ,
  \246(160) ,
  \148(851) ,
  \257(171) ,
  \290(704) ,
  \411(264) ,
  \280(850) ,
  \237(309) ,
  \173(389) ,
  \179(118) ,
  \308(1425) ,
  \268(178) ,
  \221(305) ,
  \158(349) ,
  \279(189) ,
  \214(151) ,
  \331(1401) ,
  \241(155) ,
  \190(127) ,
  \174(115) ,
  \305(702) ,
  \185(124) ,
  \263(173) ,
  \196(133) ,
  \171(621) ,
  \210(147) ,
  \169(114) ,
  \205(142) ,
  \252(166) ,
  \227(1179) ,
  \274(184) ,
  \166(625) ,
  \223(413) ,
  \247(161) ,
  \238(304) ,
  \286(696) ,
  \395(1392) ;
wire
  \2778(711) ,
  \1681(380) ,
  \1679(479) ,
  \2501(357) ,
  \1014(877) ,
  \539(1042) ,
  \600(891) ,
  \2262(689) ,
  \1243(828) ,
  \1361(1038) ,
  \1586(839) ,
  \822(497) ,
  \2422(783) ,
  \2562(727) ,
  \695(1102) ,
  \1891(1088) ,
  \616(1146) ,
  \2662(679) ,
  \1583(916) ,
  \2414(1234) ,
  \2642(603) ,
  \1932(983) ,
  \216(333) ,
  \1235(733) ,
  \537(945) ,
  \2719(1190) ,
  \825(399) ,
  \2646(675) ,
  \699(1030) ,
  \1538(580) ,
  \1984(271) ,
  \1208(1412) ,
  \900(1270) ,
  \2130(875) ,
  \643(1379) ,
  \2035(519) ,
  \2746(717) ,
  \1546(729) ,
  \1621(1055) ,
  \1225(660) ,
  \2032(634) ,
  \2122(774) ,
  \2549(962) ,
  \1238(1416) ,
  \1809(662) ,
  \2184(881) ,
  \2762(716) ,
  \1447(475) ,
  \2321(1320) ,
  \1740(535) ,
  \1979(273) ,
  \462(802) ,
  \679(1210) ,
  \1174(1327) ,
  \2161(707) ,
  \1172(1295) ,
  \671(1202) ,
  \570(890) ,
  \682(1367) ,
  \1110(1211) ,
  \1567(920) ,
  \646(1254) ,
  \2749(437) ,
  \1716(407) ,
  \2283(1156) ,
  \2665(582) ,
  \1551(1062) ,
  \1938(973) ,
  \1444(384) ,
  \1767(925) ,
  \731(1013) ,
  \1806(587) ,
  \1746(528) ,
  \2278(1130) ,
  \989(1409) ,
  \1763(857) ,
  \1781(574) ,
  \1695(482) ,
  \705(942) ,
  \1089(1423) ,
  \1600(981) ,
  \1701(556) ,
  \2177(790) ,
  \2282(1191) ,
  \2512(355) ,
  \917(1268) ,
  \982(1394) ,
  \1558(1053) ,
  \675(1060) ,
  \1167(1371) ,
  \466(667) ,
  \1549(963) ,
  \1337(898) ,
  \828(499) ,
  \2607(358) ,
  \1143(1266) ,
  \2051(738) ,
  \2214(1025) ,
  \2495(270) ,
  \2606(812) ,
  \1484(329) ,
  \2363(1159) ,
  \1589(746) ,
  \2054(970) ,
  \1822(820) ,
  \2479(278) ,
  \2140(943) ,
  \2546(743) ,
  \1430(336) ,
  \2622(811) ,
  \1333(571) ,
  \2765(433) ,
  \973(1361) ,
  \1623(998) ,
  \1049(622) ,
  \1179(1294) ,
  \2176(776) ,
  \1536(665) ,
  \2528(550) ,
  \2733(961) ,
  \560(295) ,
  \1517(447) ,
  \1743(642) ,
  \702(1176) ,
  \1547(652) ,
  \1369(1004) ,
  \1690(463) ,
  \714(1105) ,
  \2449(238) ,
  \1197(1385) ,
  \2493(361) ,
  \505(1067) ,
  \468(797) ,
  \2038(635) ,
  \2477(369) ,
  \1528(578) ,
  \1556(1111) ,
  \2623(354) ,
  \1771(766) ,
  \723(863) ,
  \2433(242) ,
  \2362(1194) ,
  \1529(592) ,
  \1498(417) ,
  \1570(843) ,
  \908(1248) ,
  \2469(458) ,
  \1870(982) ,
  \610(1024) ,
  \510(1014) ,
  \2154(631) ,
  \1939(1229) ,
  \1240(1417) ,
  \1313(503) ,
  \1550(901) ,
  \486(312) ,
  \2025(522) ,
  \983(1389) ,
  \2707(428) ,
  \2147(888) ,
  \1707(558) ,
  \152(599) ,
  \1027(1407) ,
  \2061(906) ,
  \2717(1018) ,
  \1196(1355) ,
  \916(1252) ,
  \995(798) ,
  \2060(829) ,
  \1698(563) ,
  \1091(1045) ,
  \1626(1119) ,
  \1377(997) ,
  \1974(275) ,
  \522(1171) ,
  \2270(1134) ,
  \2730(546) ,
  \964(1344) ,
  \1898(958) ,
  \2160(778) ,
  \1028(617) ,
  \2302(1174) ,
  \2215(1009) ,
  \175(710) ,
  \2113(795) ,
  \2207(759) ,
  \994(412) ,
  \1876(972) ,
  \1749(644) ,
  \534(1100) ,
  \2159(892) ,
  \2353(1243) ,
  \2273(1215) ,
  \1969(277) ,
  \827(510) ,
  \1186(1360) ,
  \1918(1052) ,
  \1247(1418) ,
  \665(1260) ,
  \1473(545) ,
  \625(1076) ,
  \1099(1259) ,
  \1816(1127) ,
  \641(1365) ,
  \1592(987) ,
  \1513(593) ,
  \2502(359) ,
  \1601(960) ,
  \580(1023) ,
  \1588(990) ,
  \1442(483) ,
  \147(600) ,
  \1453(468) ,
  \1912(959) ,
  \1133(1131) ,
  \1887(1086) ,
  \553(554) ,
  \711(946) ,
  \1311(493) ,
  \1947(1091) ,
  \1088(1421) ,
  \2525(549) ,
  \2599(360) ,
  \1355(957) ,
  \2216(1065) ,
  \729(856) ,
  \2505(266) ,
  \2258(870) ,
  \2419(1182) ,
  \742(951) ,
  \1518(551) ,
  \558(400) ,
  \2490(276) ,
  \926(1269) ,
  \1696(473) ,
  \2417(1328) ,
  \2266(775) ,
  \2313(1223) ,
  \1116(1376) ,
  \1385(283) ,
  \1893(410) ,
  \2598(813) ,
  \2518(418) ,
  \707(1043) ,
  \2167(796) ,
  \2393(1226) ,
  \1941(1228) ,
  \1060(626) ,
  \2299(1164) ,
  \664(1312) ,
  \1928(989) ,
  \1598(836) ,
  \2727(899) ,
  \1693(382) ,
  \1907(954) ,
  \1579(917) ,
  \1477(421) ,
  \2334(784) ,
  \2638(602) ,
  \969(1359) ,
  \2567(368) ,
  \2044(833) ,
  \2041(911) ,
  \1951(1089) ,
  \2339(1184) ,
  \1736(536) ,
  \599(865) ,
  \1525(540) ,
  \737(1015) ,
  \883(668) ,
  \1314(395) ,
  \834(491) ,
  \2047(740) ,
  \2426(872) ,
  \502(855) ,
  \1617(1057) ,
  \1537(654) ,
  \2382(1154) ,
  \1561(754) ,
  \1043(693) ,
  \2242(1187) ,
  \2566(819) ,
  \2137(882) ,
  \885(596) ,
  \1572(1002) ,
  \2690(348) ,
  \2366(1132) ,
  \1619(1001) ,
  \676(1006) ,
  \1881(1095) ,
  \2134(787) ,
  \979(1352) ,
  \1655(243) ,
  \2655(613) ,
  \2634(555) ,
  \1320(516) ,
  \2582(818) ,
  \2028(638) ,
  \1092(1106) ,
  \1820(739) ,
  \624(1143) ,
  \1595(913) ,
  \648(1366) ,
  \1155(1167) ,
  \1165(1356) ,
  \2583(364) ,
  \2259(1186) ,
  \632(1198) ,
  \554(581) ,
  \1114(1309) ,
  \2675(261) ,
  \1710(316) ,
  \1680(470) ,
  \1817(1066) ,
  \1795(547) ,
  \1461(559) ,
  \2718(965) ,
  \2121(869) ,
  \1728(406) ,
  \837(393) ,
  \2315(1281) ,
  \2378(1196) ,
  \1850(956) ,
  \1218(583) ,
  \1761(763) ,
  \2031(524) ,
  \949(1369) ,
  \2129(786) ,
  \1485(330) ,
  \2734(584) ,
  \1964(279) ,
  \1329(569) ,
  \2494(363) ,
  \584(1074) ,
  \2725(1247) ,
  \1739(647) ,
  \1206(1410) ,
  \1195(1350) ,
  \1879(1224) ,
  \508(858) ,
  \1793(432) ,
  \1066(627) ,
  \2148(884) ,
  \1108(1007) ,
  \1094(903) ,
  \772(297) ,
  \2464(287) ,
  \889(670) ,
  \2434(241) ,
  \2206(1149) ,
  \990(1402) ,
  \2637(683) ,
  \2402(1236) ,
  \2110(685) ,
  \2626(718) ,
  \1456(387) ,
  \1068(701) ,
  \1866(988) ,
  \2682(233) ,
  \2629(440) ,
  \1842(1037) ,
  \1418(244) ,
  \688(1381) ,
  \854(566) ,
  \1753(674) ,
  \2379(1161) ,
  \1686(462) ,
  \629(1199) ,
  \2691(252) ,
  \640(1246) ,
  \1382(1116) ,
  \2286(1138) ,
  \925(1265) ,
  \2708(427) ,
  \838(564) ,
  \562(672) ,
  \1207(1403) ,
  \684(1258) ,
  \821(390) ,
  \886(757) ,
  \2195(948) ,
  \1829(966) ,
  \2686(258) ,
  \2653(678) ,
  \2467(371) ,
  \1845(953) ,
  \528(1172) ,
  \1443(474) ,
  \2331(1181) ,
  \2291(1157) ,
  \2459(325) ,
  \1566(844) ,
  \1721(315) ,
  \2735(352) ,
  \962(1314) ,
  \1582(840) ,
  \1181(1261) ,
  \637(1245) ,
  \1557(1093) ,
  \2007(405) ,
  \1563(921) ,
  \1309(502) ,
  \1109(1123) ,
  \2227(1308) ,
  \735(859) ,
  \1691(481) ,
  \1205(1388) ,
  \1126(1249) ,
  \2398(1177) ,
  \680(1363) ,
  \1232(659) ,
  \683(1310) ,
  \1325(505) ,
  \2290(1195) ,
  \2057(907) ,
  \1532(666) ,
  \634(1256) ,
  \638(1188) ,
  \1175(1372) ,
  \2070(260) ,
  \2037(523) ,
  \2674(734) ,
  \1545(822) ,
  \2289(1213) ,
  \2610(725) ,
  \2164(686) ,
  \157(259) ,
  \1245(826) ,
  \987(1404) ,
  \655(319) ,
  \2450(237) ,
  \1959(281) ,
  \1467(561) ,
  \2369(1216) ,
  \1542(731) ,
  \2050(971) ,
  \852(619) ,
  \2234(1263) ,
  \1585(747) ,
  \2513(441) ,
  \1758(924) ,
  \2699(248) ,
  \1112(1339) ,
  \1490(542) ,
  \601(930) ,
  \154(964) ,
  \1624(1120) ,
  \2251(1183) ,
  \2613(444) ,
  \981(1377) ,
  \2470(456) ,
  \2018(404) ,
  \1934(980) ,
  \2099(249) ,
  \1025(1399) ,
  \1213(585) ,
  \2370(1192) ,
  \897(755) ,
  \2175(871) ,
  \1861(1049) ,
  \999(895) ,
  \1085(1408) ,
  \1742(530) ,
  \2141(793) ,
  \2705(339) ,
  \824(508) ,
  \2550(835) ,
  \1754(854) ,
  \967(1204) ,
  \547(415) ,
  \1449(467) ,
  \2034(633) ,
  \1307(492) ,
  \633(1142) ,
  \1087(1275) ,
  \1524(579) ,
  \456(709) ,
  \1164(1169) ,
  \2766(808) ,
  \2371(1160) ,
  \687(1357) ,
  \650(1380) ,
  \1118(1274) ,
  \1182(1343) ,
  \2639(605) ,
  \2551(372) ,
  \972(1347) ,
  \2565(455) ,
  \1317(459) ,
  \1475(331) ,
  \2541(902) ,
  \882(317) ,
  \2581(452) ,
  \1872(979) ,
  \2759(345) ,
  \819(509) ,
  \2775(341) ,
  \2524(576) ,
  \2310(1173) ,
  \922(1137) ,
  \1689(381) ,
  \1189(1348) ,
  \1568(1005) ,
  \609(867) ,
  \1454(486) ,
  \1323(496) ,
  \2390(1178) ,
  \2782(804) ,
  \2138(880) ,
  \1856(1051) ,
  \1316(515) ,
  \1072(628) ,
  \2158(708) ,
  \1335(572) ,
  \571(929) ,
  \2673(769) ,
  \2205(1147) ,
  \2056(830) ,
  \823(518) ,
  \2318(1231) ,
  \1106(1201) ,
  \2185(940) ,
  \2281(1212) ,
  \1745(641) ,
  \1762(764) ,
  \2225(1148) ,
  \2361(1219) ,
  \552(460) ,
  \613(1078) ,
  \1371(1056) ,
  \1794(430) ,
  \1643(337) ,
  \605(1022) ,
  \592(760) ,
  \1227(681) ,
  \1885(1087) ,
  \1573(751) ,
  \1925(992) ,
  \988(1387) ,
  \1273(377) ,
  \2338(873) ,
  \1828(1048) ,
  \2750(809) ,
  \2535(825) ,
  \1074(703) ,
  \2401(1227) ,
  \1748(534) ,
  \473(1420) ,
  \1826(1299) ,
  \2586(722) ,
  \1584(993) ,
  \1560(1221) ,
  \2076(257) ,
  \579(866) ,
  \1156(1297) ,
  \896(846) ,
  \807(375) ,
  \1326(398) ,
  \1945(1096) ,
  \1117(1251) ,
  \1035(618) ,
  \1864(1112) ,
  \2027(525) ,
  \1457(425) ,
  \826(489) ,
  \575(1021) ,
  \2478(234) ,
  \1692(472) ,
  \2650(606) ,
  \690(1393) ,
  \642(1345) ,
  \947(1353) ,
  \2716(928) ,
  \1148(1323) ,
  \2654(677) ,
  \1801(1017) ,
  \2468(373) ,
  \2347(1185) ,
  \1368(1058) ,
  \525(1029) ,
  \1146(1298) ,
  \743(800) ,
  \1594(837) ,
  \2403(1285) ,
  \971(1336) ,
  \1078(629) ,
  \1575(918) ,
  \2267(1158) ,
  \2062(968) ,
  \1194(1383) ,
  \2040(834) ,
  \1389(610) ,
  \948(1319) ,
  \2059(736) ,
  \1555(1064) ,
  \2503(445) ,
  \1256(401) ,
  \701(1103) ,
  \492(1035) ,
  \588(936) ,
  \2697(342) ,
  \1553(1110) ,
  \1509(552) ,
  \1310(394) ,
  \2043(741) ,
  \954(1289) ,
  \1521(541) ,
  \2210(933) ,
  \881(408) ,
  \1158(1324) ,
  \2533(664) ,
  \830(490) ,
  \2554(724) ,
  \2190(792) ,
  \1394(246) ,
  \1250(604) ,
  \1188(1337) ,
  \2323(1282) ,
  \1827(1238) ,
  \2726(1107) ,
  \2570(723) ,
  \2715(904) ,
  \2224(1080) ,
  \2374(1140) ,
  \639(1126) ,
  \2114(771) ,
  \2103(247) ,
  \2024(636) ,
  \1818(1011) ,
  \2738(714) ,
  \1591(914) ,
  \1378(1121) ,
  \1578(841) ,
  \2157(777) ,
  \1127(1271) ,
  \1507(453) ,
  \898(756) ,
  \2706(340) ,
  \1687(480) ,
  \725(1020) ,
  \1173(1354) ,
  \1863(991) ,
  \1119(1304) ,
  \833(392) ,
  \2614(817) ,
  \490(886) ,
  \1877(1225) ,
  \1544(651) ,
  \2123(697) ,
  \1261(296) ,
  \2754(713) ,
  \708(1104) ,
  \748(411) ,
  \1406(338) ,
  \2168(772) ,
  \2709(827) ,
  \1500(538) ,
  \2514(439) ,
  \937(1163) ,
  \2487(274) ,
  \980(1384) ,
  \2387(1168) ,
  \1920(995) ,
  \1147(1283) ,
  \2663(767) ,
  \2770(712) ,
  \2204(1079) ,
  \2712(861) ,
  \649(1346) ,
  \1682(469) ,
  \968(1333) ,
  \155(967) ,
  \1455(477) ,
  \1495(419) ,
  \795(294) ,
  \2757(435) ,
  \1784(436) ,
  \957(1370) ,
  \2615(356) ,
  \1786(548) ,
  \1180(1313) ,
  \749(801) ,
  \769(878) ,
  \2773(431) ,
  \1016(938) ,
  \1776(323) ,
  \2065(715) ,
  \2322(1290) ,
  \732(1068) ,
  \1541(577) ,
  \1380(1118) ,
  \2046(974) ,
  \978(1349) ,
  \1752(762) ,
  \2307(1166) ,
  \1735(645) ,
  \1452(386) ,
  \1476(332) ,
  \1113(1368) ,
  \2485(365) ,
  \504(1012) ,
  \2337(1239) ,
  \2630(810) ,
  \1057(624) ,
  \1157(1284) ,
  \2241(770) ,
  \1858(994) ,
  \1344(286) ,
  \2471(282) ,
  \487(403) ,
  \887(597) ,
  \1107(1061) ,
  \940(1318) ,
  \1738(531) ,
  \551(544) ,
  \2538(730) ,
  \930(1317) ,
  \1704(557) ,
  \1751(643) ,
  \1140(1139) ,
  \1199(1395) ,
  \1080(705) ,
  \2082(255) ,
  \2460(326) ,
  \2498(272) ,
  \963(1262) ,
  \2741(438) ,
  \2457(236) ,
  \1193(1374) ,
  \2186(944) ,
  \1562(845) ,
  \767(937) ,
  \1319(495) ,
  \1597(744) ,
  \1825(821) ,
  \977(1382) ,
  \2297(1214) ,
  \2001(314) ,
  \2441(240) ,
  \927(1315) ,
  \2033(520) ,
  \516(616) ,
  \674(1200) ,
  \894(533) ,
  \1321(504) ,
  \836(501) ,
  \2053(908) ,
  \608(932) ,
  \2671(658) ,
  \1607(1040) ,
  \2298(1208) ,
  \2377(1217) ,
  \1142(1153) ,
  \1836(955) ,
  \569(864) ,
  \820(498) ,
  \1921(1115) ,
  \1096(905) ,
  \1930(986) ,
  \2482(280) ,
  \1460(335) ,
  \1554(1063) ,
  \1100(1341) ,
  \1041(620) ,
  \144(601) ,
  \681(1340) ,
  \1614(1059) ,
  \696(1175) ,
  \2226(1150) ,
  \2257(1241) ,
  \1581(748) ,
  \1559(1109) ,
  \738(1071) ,
  \2668(614) ,
  \2203(1081) ,
  \546(322) ,
  \2223(1082) ,
  \2012(313) ,
  \970(1332) ,
  \1569(752) ,
  \1955(320) ,
  \496(862) ,
  \511(1070) ,
  \578(931) ,
  \901(1303) ,
  \1445(466) ,
  \1814(1069) ,
  \2522(539) ,
  \1868(985) ,
  \1450(485) ,
  \2115(780) ,
  \1936(976) ,
  \1481(543) ,
  \2172(690) ,
  \2504(443) ,
  \2030(637) ,
  \2088(253) ,
  \1187(1334) ,
  \835(512) ,
  \1254(308) ,
  \2523(653) ,
  \1128(1302) ,
  \1228(735) ,
  \1504(575) ,
  \946(1165) ,
  \1552(978) ,
  \1685(388) ,
  \1458(426) ,
  \1688(471) ,
  \1234(657) ,
  \621(1075) ,
  \2515(553) ,
  \2698(344) ,
  \2534(663) ,
  \1744(529) ,
  \1296(374) ,
  \2702(250) ,
  \2169(782) ,
  \1018(879) ,
  \540(1101) ,
  \2200(1031) ,
  \2306(1233) ,
  \2220(1032) ,
  \1741(646) ,
  \647(1307) ,
  \2131(789) ,
  \2058(969) ,
  \2326(1230) ,
  \[100] ,
  \1312(514) ,
  \918(1305) ,
  \2149(947) ,
  \628(1144) ,
  \1098(1311) ,
  \[102] ,
  \2052(831) ,
  \1508(451) ,
  \2126(785) ,
  \2521(595) ,
  \[103] ,
  \1201(1398) ,
  \976(1373) ,
  \2531(589) ,
  \1204(1405) ,
  \[104] ,
  \693(1028) ,
  \1331(570) ,
  \596(853) ,
  \[105] ,
  \2575(366) ,
  \1104(1203) ,
  \2461(285) ,
  \[106] ,
  \2558(816) ,
  \631(1255) ,
  \1580(996) ,
  \[107] ,
  \907(1133) ,
  \493(1083) ,
  \[108] ,
  \899(1250) ,
  \[109] ,
  \2508(268) ,
  \2230(1206) ,
  \891(669) ,
  \1184(1205) ,
  \2193(889) ,
  \2406(1235) ,
  \1999(265) ,
  \1051(695) ,
  \2039(742) ,
  \893(598) ,
  \928(1292) ,
  \2197(1033) ,
  \1953(1092) ,
  \[110] ,
  \713(1044) ,
  \1943(1097) ,
  \829(391) ,
  \1539(732) ,
  \938(1291) ,
  \2118(688) ,
  \1790(588) ,
  \1587(915) ,
  \2532(590) ,
  \2036(632) ,
  \2664(768) ,
  \685(1375) ,
  \498(1019) ,
  \521(1098) ,
  \635(1189) ,
  \1823(728) ,
  \2458(235) ,
  \471(1419) ,
  \2591(362) ,
  \2217(1034) ,
  \2543(900) ,
  \1115(1257) ,
  \2213(852) ,
  \1448(385) ,
  \2395(1170) ,
  \1493(327) ,
  \1322(397) ,
  \720(1084) ,
  \2574(815) ,
  \1819(1128) ,
  \984(1397) ,
  \1785(434) ,
  \1615(1003) ,
  \1257(893) ,
  \884(1386) ,
  \2233(1338) ,
  \2350(687) ,
  \2023(526) ,
  \2151(691) ,
  \2590(814) ,
  \2658(611) ,
  \2683(256) ,
  \[122] ,
  \2342(779) ,
  \2418(1293) ,
  \955(1351) ,
  \2722(1047) ,
  \1772(860) ,
  \2542(824) ,
  \909(1267) ,
  \1590(838) ,
  \[125] ,
  \2411(1286) ,
  \1571(919) ,
  \2055(737) ,
  \2618(719) ,
  \1166(1325) ,
  \1062(699) ,
  \[127] ,
  \[128] ,
  \2486(367) ,
  \480(292) ,
  \1284(293) ,
  \2275(1155) ,
  \1830(1108) ,
  \1874(975) ,
  \1678(461) ,
  \1747(640) ,
  \620(1145) ,
  \1859(1114) ,
  \1798(927) ,
  \1631(245) ,
  \1135(1272) ,
  \2631(615) ,
  \630(1141) ,
  \1006(799) ,
  \2274(1193) ,
  \677(1122) ,
  \956(1321) ,
  \[130] ,
  \1683(487) ,
  \910(1301) ,
  \1813(661) ,
  \[131] ,
  \2661(680) ,
  \2645(676) ,
  \1031(630) ,
  \1499(324) ,
  \533(1041) ,
  \1694(464) ,
  \846(565) ,
  \1464(560) ,
  \2094(251) ,
  \2743(350) ,
  \[137] ,
  \1775(416) ,
  \1824(650) ,
  \929(1279) ,
  \1574(842) ,
  \[139] ,
  \784(378) ,
  \2559(370) ,
  \2029(521) ,
  \1994(267) ,
  \2049(909) ,
  \1111(1364) ,
  \753(896) ,
  \2196(950) ,
  \939(1280) ,
  \875(290) ,
  \2605(446) ,
  \2602(720) ,
  \1200(1390) ,
  \2589(450) ,
  \857(567) ,
  \1459(424) ,
  \1093(1220) ,
  \2442(239) ,
  \2183(883) ,
  \1810(586) ,
  \2425(1240) ,
  \1540(655) ,
  \1750(527) ,
  \2180(788) ,
  \1012(935) ,
  \2694(254) ,
  \1005(952) ,
  \645(1197) ,
  \1451(476) ,
  \2355(1162) ,
  \2243(1300) ,
  \2672(682) ,
  \1543(750) ,
  \2386(1209) ,
  \1577(749) ,
  \1777(537) ,
  \1923(1050) ,
  \765(876) ,
  \895(1396) ,
  \1989(269) ,
  \258(321) ,
  \1628(1117) ,
  \2557(457) ,
  \2345(1242) ,
  \717(887) ,
  \1239(1415) ,
  \1831(409) ,
  \2621(442) ,
  \2042(977) ,
  \1134(1253) ,
  \2511(353) ,
  \686(1329) ,
  \2647(608) ,
  \2346(868) ,
  \2139(939) ,
  \146(758) ,
  \1548(823) ,
  \2026(639) ,
  \2758(806) ,
  \1734(532) ,
  \2194(885) ,
  \1351(284) ,
  \1446(484) ,
  \2410(1296) ,
  \658(318) ,
  \1315(494) ,
  \841(573) ,
  \[84] ,
  \1145(1316) ,
  \1373(1000) ,
  \1593(745) ,
  \[85] ,
  \2385(1218) ,
  \1533(591) ,
  \[86] ,
  \617(1077) ,
  \1125(1135) ,
  \[87] ,
  \[88] ,
  \1486(420) ,
  \1251(310) ,
  \[89] ,
  \2573(454) ,
  \832(500) ,
  \763(934) ,
  \1949(1090) ,
  \726(1073) ,
  \1387(594) ,
  \1327(568) ,
  \187(673) ,
  \1737(648) ,
  \719(1036) ,
  \1516(449) ,
  \636(1125) ,
  \2187(794) ,
  \1596(984) ,
  \2235(684) ,
  \2246(1207) ,
  \[90] ,
  \2294(1152) ,
  \1198(1378) ,
  \[91] ,
  \1904(1039) ,
  \2681(351) ,
  \1375(1054) ,
  \961(1288) ,
  \[92] ,
  \2767(343) ,
  \1667(334) ,
  \2409(1326) ,
  \2774(805) ,
  \[93] ,
  \1889(1085) ,
  \2265(1244) ,
  \1308(513) ,
  \2250(1264) ,
  \2107(706) ,
  \531(941) ,
  \1697(383) ,
  \[95] ,
  \1441(465) ,
  \589(1026) ,
  \[96] ,
  \[97] ,
  \2144(791) ,
  \527(1099) ,
  \[98] ,
  \644(1391) ,
  \2329(1322) ,
  \2578(726) ,
  \2048(832) ,
  \924(1151) ,
  \2045(910) ,
  \499(1072) ,
  \1144(1273) ,
  \2358(1136) ,
  \2238(1124) ,
  \1576(999) ,
  \2249(1331) ,
  \1494(328) ,
  \1815(1010) ,
  \2305(1222) ,
  \1564(1008) ,
  \475(897) ,
  \991(1411) ,
  \1565(753) ,
  \519(1027) ,
  \1770(765) ,
  \1802(926) ,
  \1805(1016) ,
  \831(511) ,
  \1185(1335) ,
  \2742(807) ,
  \1926(1113) ,
  \2254(781) ,
  \1258(894) ,
  \1221(1413) ,
  \1253(402) ,
  \1684(478) ,
  \2751(347) ,
  \2330(1287) ,
  \550(422) ,
  \1470(562) ,
  \1324(517) ,
  \1599(912) ,
  \654(300) ,
  \2314(1232) ,
  \2781(429) ,
  \2150(949) ,
  \1883(1094) ,
  \865(291) ,
  \2594(721) ,
  \666(1342) ,
  \2597(448) ,
  \587(874) ,
  \1318(396) ,
  \143(1330) ,
  \1821(649) ,
  \2394(1237) ,
  \818(488) ,
  \1190(1362) ,
  \2689(346) ,
  \2354(773) ,
  \1136(1306) ,
  \915(1129) ;
assign
  \2778(711)  = \2036(632)  | \2035(519) ,
  \1681(380)  = \1655(243)  & (\1631(245)  & \118(93) ),
  \269(179)  = \IN-269(179) ,
  \1679(479)  = \1667(334)  & (\1631(245)  & \106(83) ),
  \215(152)  = \IN-215(152) ,
  \2501(357)  = ~\2495(270) ,
  \1014(877)  = \995(798)  & \1057(624) ,
  \539(1042)  = \748(411)  & \537(945) ,
  \600(891)  = ~\2168(772)  | ~\2161(707) ,
  \2262(689)  = \1035(618) ,
  \1243(828)  = ~\1228(735) ,
  \1361(1038)  = ~\1355(957) ,
  \1586(839)  = ~\2606(812)  | ~\2599(360) ,
  \822(497)  = \807(375)  & (\784(378)  & \81(62) ),
  \2422(783)  = \1051(695) ,
  \2562(727)  = \1737(648)  | \1736(536) ,
  \695(1102)  = \994(412)  & \693(1028) ,
  \1891(1088)  = \1845(953)  & \1876(972) ,
  \616(1146)  = ~\613(1078) ,
  \2662(679)  = ~\2658(611) ,
  \1583(916)  = ~\1582(840)  | ~\1581(748) ,
  \2414(1234)  = \696(1175) ,
  \2642(603)  = \1701(556) ,
  \1932(983)  = \1912(959)  & \1989(269) ,
  \216(333)  = \1955(320)  & \2106(222) ,
  \1235(733)  = \1234(657)  | \1232(659) ,
  \156(1046)  = \[125] ,
  \537(945)  = \753(896)  & \1072(628) ,
  \2719(1190)  = ~\1816(1127)  | ~\1819(1128) ,
  \397(1406)  = \1025(1399) ,
  \825(399)  = \795(294)  & (\772(297)  & \68(51) ),
  \2646(675)  = ~\2642(603) ,
  \699(1030)  = \1018(879)  | \1016(938) ,
  \1538(580)  = \1521(541)  & (\1477(421)  & \1486(420) ),
  \1984(271)  = ~\1981(208) ,
  \1208(1412)  = \1207(1403)  | \1206(1410) ,
  \900(1270)  = ~\2274(1193)  | ~\2267(1158) ,
  \2130(875)  = ~\2126(785) ,
  \643(1379)  = ~\642(1345)  | ~\641(1365) ,
  \2035(519)  = \2018(404)  & \35(26) ,
  \2746(717)  = \2028(638)  | \2027(525) ,
  \1546(729)  = \1536(665)  & (\1513(593)  & \1500(538) ),
  \1621(1055)  = \1607(1040)  & \2082(255) ,
  \1225(660)  = \1213(585)  & \2099(249) ,
  \2032(634)  = \2012(313)  & \1461(559) ,
  \2122(774)  = ~\2118(688) ,
  \2549(962)  = ~\2543(900) ,
  \1238(1416)  = \1221(1413)  & \1208(1412) ,
  \1809(662)  = ~\1806(587) ,
  \2184(881)  = ~\2180(788) ,
  \2762(716)  = \2032(634)  | \2031(524) ,
  \1447(475)  = \1418(244)  & (\1406(338)  & \125(98) ),
  \2321(1320)  = ~\2315(1281) ,
  \1740(535)  = \1716(407)  & \5(4) ,
  \1979(273)  = ~\1976(207) ,
  \462(802)  = ~\456(709) ,
  \679(1210)  = \1031(630)  & \677(1122) ,
  \1174(1327)  = ~\2418(1293)  | ~\2411(1286) ,
  \2161(707)  = \1031(630) ,
  \1172(1295)  = \702(1176)  & \1941(1228) ,
  \671(1202)  = \1043(693)  & \1380(1118) ,
  \570(890)  = ~\2114(771)  | ~\2107(706) ,
  \682(1367)  = \679(1210)  & (\666(1342)  & \681(1340) ),
  \1110(1211)  = \1031(630)  & \1109(1123) ,
  \180(119)  = \IN-180(119) ,
  \145(1358)  = \[131] ,
  \1567(920)  = ~\1566(844)  | ~\1565(753) ,
  \646(1254)  = ~\2242(1187)  | ~\2235(684) ,
  \2749(437)  = ~\2743(350) ,
  \1716(407)  = ~\1710(316) ,
  \2283(1156)  = \1887(1086) ,
  \2665(582)  = \1473(545) ,
  \1551(1062)  = ~\2549(962)  | ~\2546(743) ,
  \1938(973)  = \1912(959)  & \2070(260) ,
  \1444(384)  = \1418(244)  & (\1394(246)  & \114(89) ),
  \1767(925)  = ~\1763(857) ,
  \731(1013)  = \1005(952)  & \729(856) ,
  \1806(587)  = \1795(547) ,
  \1746(528)  = \1728(406)  & \23(16) ,
  \191(128)  = \IN-191(128) ,
  \2278(1130)  = \505(1067) ,
  \989(1409)  = \987(1404)  & \973(1361) ,
  \1763(857)  = ~\1762(764)  | ~\1761(763) ,
  \1781(574)  = ~\1777(537) ,
  \1695(482)  = \1667(334)  & (\1631(245)  & \103(80) ),
  \705(942)  = \999(895)  & \1066(627) ,
  \1089(1423)  = \554(581)  & (\1088(1421)  & \1085(1408) ),
  \1600(981)  = ~\1599(912) ,
  \1701(556)  = \1689(381)  | (\1688(471)  | (\1687(480)  | \1686(462) )),
  \2177(790)  = \1068(701) ,
  \200(137)  = \IN-200(137) ,
  \186(125)  = \IN-186(125) ,
  \2282(1191)  = ~\2278(1130) ,
  \2512(355)  = ~\2508(268) ,
  \917(1268)  = ~\2290(1195)  | ~\2283(1156) ,
  \982(1394)  = \981(1377)  | (\980(1384)  | (\979(1352)  | (\978(1349)  | \937(1163) ))),
  \1558(1053)  = \2042(977)  & (\2046(974)  & (\2050(971)  & (\2054(970)  & \2058(969) ))),
  \675(1060)  = \1361(1038)  & \1999(265) ,
  \1167(1371)  = ~\1166(1325)  | ~\1165(1356) ,
  \466(667)  = ~\1387(594) ,
  \1549(963)  = ~\2541(902)  | ~\2538(730) ,
  \1337(898)  = \462(802) ,
  \828(499)  = \795(294)  & (\784(378)  & \66(49) ),
  \197(134)  = \IN-197(134) ,
  \2607(358)  = \1984(271) ,
  \1143(1266)  = ~\2385(1218)  | ~\2382(1154) ,
  \242(156)  = \IN-242(156) ,
  \2051(738)  = ~\2765(433)  | ~\2762(716) ,
  \264(174)  = \IN-264(174) ,
  \2214(1025)  = ~\2210(933) ,
  \2495(270)  = \1986(209) ,
  \2606(812)  = ~\2602(720) ,
  \1484(329)  = ~\2441(240)  | ~\2438(226) ,
  \2363(1159)  = \1951(1089) ,
  \1589(746)  = ~\2613(444)  | ~\2610(725) ,
  \2054(970)  = ~\2053(908) ,
  \1822(820)  = ~\1821(649)  & ~\1820(739) ,
  \2479(278)  = \1966(205) ,
  \2140(943)  = ~\2138(880)  | ~\2131(789) ,
  \211(148)  = \IN-211(148) ,
  \2546(743)  = ~\2534(663)  | ~\2533(664) ,
  \206(143)  = \IN-206(143) ,
  \1430(336)  = ~\1418(244) ,
  \2622(811)  = ~\2618(719) ,
  \253(167)  = \IN-253(167) ,
  \1333(571)  = \1322(397)  | (\1321(504)  | (\1320(516)  | \1319(495) )),
  \275(185)  = \IN-275(185) ,
  \2765(433)  = ~\2759(345) ,
  \973(1361)  = \972(1347)  | (\971(1336)  | (\970(1332)  | \907(1133) )),
  \1623(998)  = \1601(960)  & \1964(279) ,
  \1049(622)  = \857(567) ,
  \1179(1294)  = \696(1175)  & \1939(1229) ,
  \2176(776)  = ~\2172(690) ,
  \248(162)  = \IN-248(162) ,
  \1536(665)  = ~\1533(591) ,
  \2528(550)  = ~\2504(443)  | ~\2503(445) ,
  \2733(961)  = ~\2727(899) ,
  \560(295)  = ~\559(193) ,
  \1517(447)  = ~\2494(363)  | ~\2487(274) ,
  \1743(642)  = \1721(315)  & \1327(568) ,
  \702(1176)  = ~\701(1103) ,
  \1547(652)  = \1533(591)  & (\1504(575)  & \1513(593) ),
  \1369(1004)  = \1355(957)  & \1351(284) ,
  \1690(463)  = \1667(334)  & (\1643(337)  & \140(111) ),
  \714(1105)  = ~\713(1044) ,
  \2449(238)  = ~\2443(227) ,
  \1197(1385)  = \1158(1324)  & (\1179(1294)  & (\1148(1323)  & \1167(1371) )),
  \2493(361)  = ~\2487(274) ,
  \505(1067)  = ~\504(1012) ,
  \468(797)  = \466(667)  & (\1389(610)  & \40(29) ),
  \2038(635)  = \2012(313)  & \1470(562) ,
  \2477(369)  = ~\2471(282) ,
  \1528(578)  = ~\1525(540) ,
  \1556(1111)  = \1555(1064)  & \1554(1063) ,
  \311(1278)  = \1560(1221) ,
  \2623(354)  = \1994(267) ,
  \1771(766)  = ~\2654(677)  | ~\2647(608) ,
  \723(863)  = \1006(799)  & \1698(563) ,
  \2433(242)  = ~\2427(223) ,
  \2362(1194)  = ~\2358(1136) ,
  \1529(592)  = \1518(551) ,
  \367(288)  = \1083(199) ,
  \1498(417)  = ~\2477(369)  | ~\2474(231) ,
  \1570(843)  = ~\2574(815)  | ~\2567(368) ,
  \908(1248)  = ~\2281(1212)  | ~\2278(1130) ,
  \2469(458)  = ~\2467(371)  | ~\2464(287) ,
  \1870(982)  = \1850(956)  & \1989(269) ,
  \610(1024)  = ~\609(867)  | ~\608(932) ,
  \510(1014)  = \742(951)  & \508(858) ,
  \301(694)  = \1049(622) ,
  \225(1424)  = \[139] ,
  \2154(631)  = \841(573) ,
  \1939(1229)  = \1893(410)  & \1921(1115) ,
  \1240(1417)  = \1239(1415)  | \1238(1416) ,
  \1313(503)  = \1284(293)  & (\1273(377)  & \62(45) ),
  \1550(901)  = ~\2542(824)  | ~\2535(825) ,
  \486(312)  = \37(28) ,
  \2025(522)  = \2007(405)  & \32(23) ,
  \983(1389)  = \685(1375)  & \977(1382) ,
  \2707(428)  = ~\2705(339)  | ~\2702(250) ,
  \2147(888)  = ~\2141(793) ,
  \1707(558)  = \1697(383)  | (\1696(473)  | (\1695(482)  | \1694(464) )),
  \401(1276)  = \1093(1220) ,
  \152(599)  = \860(197)  & \841(573) ,
  \1027(1407)  = ~\1025(1399) ,
  \2061(906)  = ~\2060(829)  | ~\2059(736) ,
  \2717(1018)  = ~\2715(904)  | ~\2712(861) ,
  \1196(1355)  = \1172(1295)  & (\1148(1323)  & \1158(1324) ),
  \916(1252)  = ~\2289(1213)  | ~\2286(1138) ,
  \995(798)  = \456(709) ,
  \2060(829)  = ~\2782(804)  | ~\2775(341) ,
  \1698(563)  = \1685(388)  | (\1684(478)  | (\1683(487)  | \1682(469) )),
  \1091(1045)  = ~\1550(901)  | ~\1549(963) ,
  \1626(1119)  = \1619(1001)  | \1617(1057) ,
  \1377(997)  = \1355(957)  & \1964(279) ,
  \1974(275)  = ~\1971(206) ,
  \522(1171)  = ~\521(1098) ,
  \2270(1134)  = \511(1070) ,
  \2730(546)  = ~\2708(427)  | ~\2707(428) ,
  \964(1344)  = ~\963(1262)  | ~\962(1314) ,
  \1898(958)  = \1337(898) ,
  \2160(778)  = ~\2158(708)  | ~\2151(691) ,
  \1028(617)  = ~\838(564) ,
  \2302(1174)  = \540(1101) ,
  \2215(1009)  = ~\2213(852)  | ~\2210(933) ,
  \175(710)  = \554(581)  & (\36(27)  & (\483(191)  & \480(292) )),
  \2113(795)  = ~\2107(706) ,
  \2207(759)  = ~\562(672) ,
  \994(412)  = \655(319) ,
  \1876(972)  = \1850(956)  & \2070(260) ,
  \1749(644)  = \1721(315)  & \1333(571) ,
  \534(1100)  = ~\533(1041) ,
  \2159(892)  = ~\2157(777)  | ~\2154(631) ,
  \2353(1243)  = ~\2347(1185) ,
  \2273(1215)  = ~\2267(1158) ,
  \1969(277)  = ~\1966(205) ,
  \827(510)  = \807(375)  & (\772(297)  & \54(39) ),
  \1186(1360)  = ~\1185(1335) ,
  \1918(1052)  = \1904(1039)  & \2088(253) ,
  \1247(1418)  = ~\1240(1417) ,
  \665(1260)  = ~\2258(870)  | ~\2251(1183) ,
  \1473(545)  = \1460(335)  | (\1459(424)  | (\1458(426)  | \1457(425) )),
  \625(1076)  = \610(1024) ,
  \181(120)  = \IN-181(120) ,
  \1099(1259)  = ~\2346(868)  | ~\2339(1184) ,
  \1816(1127)  = ~\1815(1010)  & ~\1814(1069) ,
  \641(1365)  = ~\2233(1338)  | ~\2230(1206) ,
  \1592(987)  = ~\1591(914) ,
  \1513(593)  = ~\1509(552) ,
  \2502(359)  = ~\2498(272) ,
  \1601(960)  = \1337(898) ,
  \580(1023)  = ~\579(866)  | ~\578(931) ,
  \1588(990)  = ~\1587(915) ,
  \1442(483)  = \1430(336)  & (\1394(246)  & \102(79) ),
  \147(600)  = \860(197)  & \846(565) ,
  \1453(468)  = \1430(336)  & (\1406(338)  & \135(106) ),
  \1912(959)  = \1337(898) ,
  \1133(1131)  = \732(1068)  & \1951(1089) ,
  \391(379)  = \654(300) ,
  \1887(1086)  = \1845(953)  & \1872(979) ,
  \553(554)  = ~\552(460) ,
  \711(946)  = \999(895)  & \1072(628) ,
  \1311(493)  = \1296(374)  & (\1273(377)  & \88(67) ),
  \1947(1091)  = \1907(954)  & \1932(983) ,
  \1088(1421)  = \473(1420)  & (\1087(1275)  & \1553(1110) ),
  \2525(549)  = ~\2514(439)  | ~\2513(441) ,
  \2599(360)  = \1979(273) ,
  \1355(957)  = \475(897) ,
  \2216(1065)  = ~\2214(1025)  | ~\2207(759) ,
  \729(856)  = \1006(799)  & \1701(556) ,
  \2505(266)  = \1996(211) ,
  \2258(870)  = ~\2254(781) ,
  \2419(1182)  = \1628(1117) ,
  \742(951)  = \1257(893) ,
  \1518(551)  = ~\1517(447)  | ~\1516(449) ,
  \270(180)  = \IN-270(180) ,
  \558(400)  = \1251(310)  & \1254(308) ,
  \2490(276)  = \1971(206) ,
  \926(1269)  = ~\2298(1208)  | ~\2291(1157) ,
  \1696(473)  = \1655(243)  & (\1643(337)  & \127(100) ),
  \2417(1328)  = ~\2411(1286) ,
  \2266(775)  = ~\2262(689) ,
  \2313(1223)  = ~\2307(1166) ,
  \1116(1376)  = \1113(1368)  | (\1111(1364)  | \1104(1203) ),
  \1385(283)  = ~\1384(202) ,
  \1893(410)  = \658(318) ,
  \2598(813)  = ~\2594(721) ,
  \2518(418)  = ~\2460(326)  | ~\2459(325) ,
  \707(1043)  = \994(412)  & \705(942) ,
  \2167(796)  = ~\2161(707) ,
  \2393(1226)  = ~\2387(1168) ,
  \1941(1228)  = \1893(410)  & \1926(1113) ,
  \1060(626)  = \1329(569) ,
  \2299(1164)  = \1883(1094) ,
  \664(1312)  = ~\2257(1241)  | ~\2254(781) ,
  \1928(989)  = \1898(958)  & \1979(273) ,
  \1598(836)  = ~\2630(810)  | ~\2623(354) ,
  \2727(899)  = ~\1822(820)  | ~\1825(821) ,
  \1693(382)  = \1655(243)  & (\1631(245)  & \116(91) ),
  \1907(954)  = \1258(894) ,
  \1579(917)  = ~\1578(841)  | ~\1577(749) ,
  \1477(421)  = ~\1476(332)  | ~\1475(331) ,
  \2334(784)  = \1051(695) ,
  \2638(602)  = ~\2634(555) ,
  \969(1359)  = ~\968(1333) ,
  \2567(368)  = \1959(281) ,
  \2044(833)  = ~\2750(809)  | ~\2743(350) ,
  \2041(911)  = ~\2040(834)  | ~\2039(742) ,
  \1951(1089)  = \1907(954)  & \1936(976) ,
  \2339(1184)  = \1626(1119) ,
  \1736(536)  = \1716(407)  & \4(3) ,
  \162(612)  = \[103] ,
  \599(865)  = ~\2167(796)  | ~\2164(686) ,
  \1525(540)  = \1495(419) ,
  \737(1015)  = \1005(952)  & \735(859) ,
  \883(668)  = \875(290)  & \516(616) ,
  \1314(395)  = \1284(293)  & (\1261(296)  & \75(56) ),
  \834(491)  = \807(375)  & (\784(378)  & \90(69) ),
  \2047(740)  = ~\2757(435)  | ~\2754(713) ,
  \2426(872)  = ~\2422(783) ,
  \502(855)  = \743(800)  & \1701(556) ,
  \1617(1057)  = \1607(1040)  & \2076(257) ,
  \192(129)  = \IN-192(129) ,
  \1537(654)  = \1524(579)  & (\1486(420)  & \1481(543) ),
  \2382(1154)  = \720(1084) ,
  \1561(754)  = ~\2557(457)  | ~\2554(724) ,
  \1043(693)  = ~\1041(620) ,
  \2242(1187)  = ~\2238(1124) ,
  \2566(819)  = ~\2562(727) ,
  \2137(882)  = ~\2131(789) ,
  \885(596)  = \875(290)  & \841(573) ,
  \1572(1002)  = ~\1571(919) ,
  \350(301)  = \452(190) ,
  \2690(348)  = ~\2686(258) ,
  \2366(1132)  = \732(1068) ,
  \1619(1001)  = \1601(960)  & \1959(281) ,
  \676(1006)  = \1355(957)  & \1344(286) ,
  \1881(1095)  = \1831(409)  & \1866(988) ,
  \2134(787)  = \1062(699) ,
  \979(1352)  = \954(1289)  & (\930(1317)  & \940(1318) ),
  \1655(243)  = \2105(221) ,
  \2655(613)  = \1467(561) ,
  \2634(555)  = \1681(380)  | (\1680(470)  | (\1679(479)  | \1678(461) )),
  \1320(516)  = \1296(374)  & (\1261(296)  & \48(33) ),
  \201(138)  = \IN-201(138) ,
  \2582(818)  = ~\2578(726) ,
  \243(157)  = \IN-243(157) ,
  \2028(638)  = \2001(314)  & \1704(557) ,
  \1092(1106)  = ~\1091(1045) ,
  \265(175)  = \IN-265(175) ,
  \1820(739)  = \1809(662)  & (\1786(548)  & \1781(574) ),
  \198(135)  = \IN-198(135) ,
  \624(1143)  = ~\621(1075) ,
  \1595(913)  = ~\1594(837)  | ~\1593(745) ,
  \648(1366)  = ~\2249(1331)  | ~\2246(1207) ,
  \1155(1167)  = \714(1105)  & \1945(1096) ,
  \1165(1356)  = ~\2409(1326)  | ~\2406(1235) ,
  \212(149)  = \IN-212(149) ,
  \2583(364)  = \1969(277) ,
  \2259(1186)  = \1378(1121) ,
  \632(1198)  = \620(1145)  & (\584(1074)  & \571(929) ),
  \554(581)  = \553(554)  & \551(544) ,
  \1114(1309)  = ~\2353(1243)  | ~\2350(687) ,
  \2675(261)  = \2067(213) ,
  \1710(316)  = \16(11) ,
  \1680(470)  = \1655(243)  & (\1643(337)  & \130(103) ),
  \1817(1066)  = \1805(1016)  & (\1767(925)  & \1754(854) ),
  \1795(547)  = ~\1794(430)  | ~\1793(432) ,
  \207(144)  = \IN-207(144) ,
  \1461(559)  = \1444(384)  | (\1443(474)  | (\1442(483)  | \1441(465) )),
  \254(168)  = \IN-254(168) ,
  \2718(965)  = ~\2716(928)  | ~\2709(827) ,
  \249(163)  = \IN-249(163) ,
  \2121(869)  = ~\2115(780) ,
  \1728(406)  = ~\1721(315) ,
  \837(393)  = \795(294)  & (\772(297)  & \77(58) ),
  \2315(1281)  = \1879(1224) ,
  \2378(1196)  = ~\2374(1140) ,
  \1850(956)  = \475(897) ,
  \168(623)  = \[106] ,
  \1218(583)  = ~\1473(545)  | ~\2103(247) ,
  \1761(763)  = ~\2645(676)  | ~\2642(603) ,
  \2031(524)  = \2018(404)  & \27(20) ,
  \284(847)  = \897(755) ,
  \949(1369)  = ~\948(1319)  | ~\947(1353) ,
  \2129(786)  = ~\2123(697) ,
  \1485(330)  = ~\2442(239)  | ~\2435(225) ,
  \2734(584)  = ~\2730(546) ,
  \1964(279)  = ~\1961(204) ,
  \1329(569)  = \1314(395)  | (\1313(503)  | (\1312(514)  | \1311(493) )),
  \2494(363)  = ~\2490(276) ,
  \584(1074)  = ~\580(1023) ,
  \2725(1247)  = ~\2719(1190) ,
  \1739(647)  = \1710(316)  & \854(566) ,
  \1206(1410)  = \1204(1405)  & \1190(1362) ,
  \1195(1350)  = \1164(1169)  & \1148(1323) ,
  \150(1277)  = \[130] ,
  \1879(1224)  = \1831(409)  & \1864(1112) ,
  \508(858)  = \743(800)  & \1250(604) ,
  \1793(432)  = ~\2697(342)  | ~\2694(254) ,
  \276(186)  = \IN-276(186) ,
  \1066(627)  = \1331(570) ,
  \2148(884)  = ~\2144(791) ,
  \1108(1007)  = \1601(960)  & \1344(286) ,
  \1094(903)  = \1245(826)  & \1235(733) ,
  \772(297)  = \543(192) ,
  \2464(287)  = \1341(200) ,
  \889(670)  = \868(198)  & \1049(622) ,
  \2434(241)  = ~\2430(224) ,
  \2206(1149)  = ~\2204(1079)  | ~\2197(1033) ,
  \990(1402)  = \984(1397)  & \988(1387) ,
  \2637(683)  = ~\2631(615) ,
  \2402(1236)  = ~\2398(1177) ,
  \2110(685)  = \1028(617) ,
  \2626(718)  = \2024(636)  | \2023(526) ,
  \1456(387)  = \1418(244)  & (\1394(246)  & \111(86) ),
  \1068(701)  = ~\1066(627) ,
  \1866(988)  = \1836(955)  & \1979(273) ,
  \2682(233)  = ~\2678(232) ,
  \2629(440)  = ~\2623(354) ,
  \1842(1037)  = ~\1836(955) ,
  \1418(244)  = \2105(221) ,
  \688(1381)  = \487(403)  & \687(1357) ,
  \854(566)  = \833(392)  | (\832(500)  | (\831(511)  | \830(490) )),
  \1753(674)  = ~\2638(602)  | ~\2631(615) ,
  \2379(1161)  = \1947(1091) ,
  \1686(462)  = \1667(334)  & (\1643(337)  & \141(112) ),
  \629(1199)  = \616(1146)  & (\580(1023)  & \575(1021) ),
  \2691(252)  = \2090(217) ,
  \640(1246)  = ~\639(1126)  & ~\638(1188) ,
  \1382(1116)  = \1377(997)  | \1375(1054) ,
  \2286(1138)  = \499(1072) ,
  \925(1265)  = ~\2297(1214)  | ~\2294(1152) ,
  \2708(427)  = ~\2706(340)  | ~\2699(248) ,
  \838(564)  = \821(390)  | (\820(498)  | (\819(509)  | \818(488) )),
  \562(672)  = ~\852(619)  | ~\560(295) ,
  \1207(1403)  = \1201(1398)  & \1205(1388) ,
  \319(656)  = \554(581) ,
  \684(1258)  = ~\2266(775)  | ~\2259(1186) ,
  \821(390)  = \795(294)  & (\772(297)  & \80(61) ),
  \886(757)  = \868(198)  & \562(672) ,
  \2195(948)  = ~\2193(889)  | ~\2190(792) ,
  \1829(966)  = ~\2734(584)  | ~\2727(899) ,
  \2686(258)  = \2072(214) ,
  \2653(678)  = ~\2647(608) ,
  \2467(371)  = ~\2461(285) ,
  \1845(953)  = \1258(894) ,
  \528(1172)  = ~\527(1099) ,
  \1443(474)  = \1418(244)  & (\1406(338)  & \126(99) ),
  \2331(1181)  = \1382(1116) ,
  \2291(1157)  = \1885(1087) ,
  \2459(325)  = ~\2457(236)  | ~\2454(230) ,
  \1566(844)  = ~\2566(819)  | ~\2559(370) ,
  \1721(315)  = \16(11) ,
  \2735(352)  = \1999(265) ,
  \962(1314)  = ~\2337(1239)  | ~\2334(784) ,
  \1582(840)  = ~\2598(813)  | ~\2591(362) ,
  \1181(1261)  = ~\2426(872)  | ~\2419(1182) ,
  \637(1245)  = ~\636(1125)  & ~\635(1189) ,
  \261(506)  = \[100] ,
  \1557(1093)  = \2062(968)  & \2065(715) ,
  \299(692)  = \1041(620) ,
  \2007(405)  = ~\2001(314) ,
  \1563(921)  = ~\1562(845)  | ~\1561(754) ,
  \1309(502)  = \1284(293)  & (\1273(377)  & \63(46) ),
  \288(700)  = \1066(627) ,
  \1109(1123)  = \1108(1007)  | \1107(1061) ,
  \2227(1308)  = ~\631(1255)  | ~\634(1256) ,
  \735(859)  = \1006(799)  & \1250(604) ,
  \1691(481)  = \1667(334)  & (\1631(245)  & \104(81) ),
  \1205(1388)  = ~\1186(1360)  | ~\1193(1374) ,
  \295(1400)  = \895(1396) ,
  \1126(1249)  = ~\2369(1216)  | ~\2366(1132) ,
  \2398(1177)  = \708(1104) ,
  \680(1363)  = \674(1200)  & \666(1342) ,
  \1232(659)  = \1218(583)  & \2103(247) ,
  \683(1310)  = ~\2265(1244)  | ~\2262(689) ,
  \1325(505)  = \1284(293)  & (\1273(377)  & \60(43) ),
  \2290(1195)  = ~\2286(1138) ,
  \2057(907)  = ~\2056(830)  | ~\2055(737) ,
  \1532(666)  = ~\1529(592) ,
  \634(1256)  = ~\633(1142)  & ~\632(1198) ,
  \638(1188)  = \628(1144)  & (\605(1022)  & \592(760) ),
  \1175(1372)  = ~\1174(1327)  | ~\1173(1354) ,
  \2070(260)  = ~\2067(213) ,
  \384(262)  = \2066(212) ,
  \2037(523)  = \2018(404)  & \28(21) ,
  \2674(734)  = ~\2672(682)  | ~\2665(582) ,
  \1545(822)  = ~\1544(651)  & ~\1543(750) ,
  \2289(1213)  = ~\2283(1156) ,
  \2610(725)  = \1749(644)  | \1748(534) ,
  \2164(686)  = \1028(617) ,
  \157(259)  = \2072(214)  & (\2078(215)  & (\2084(216)  & \2090(217) )),
  \1245(826)  = ~\1235(733) ,
  \987(1404)  = ~\984(1397) ,
  \655(319)  = \8(7) ,
  \2450(237)  = ~\2446(228) ,
  \182(121)  = \IN-182(121) ,
  \1959(281)  = ~\1956(203) ,
  \1467(561)  = \1452(386)  | (\1451(476)  | (\1450(485)  | \1449(467) )),
  \2369(1216)  = ~\2363(1159) ,
  \1542(731)  = ~\1541(577)  & ~\1540(655) ,
  \2050(971)  = ~\2049(909) ,
  \852(619)  = ~\846(565) ,
  \2234(1263)  = ~\2230(1206) ,
  \193(130)  = \IN-193(130) ,
  \1585(747)  = ~\2605(446)  | ~\2602(720) ,
  \2513(441)  = ~\2511(353)  | ~\2508(268) ,
  \1758(924)  = ~\1754(854) ,
  \2699(248)  = \2100(219) ,
  \1112(1339)  = ~\1115(1257)  | ~\1114(1309) ,
  \1490(542)  = ~\1486(420) ,
  \601(930)  = ~\600(891)  | ~\599(865) ,
  \154(964)  = \1245(826)  | \1094(903) ,
  \1624(1120)  = \1615(1003)  | \1614(1059) ,
  \2251(1183)  = \1380(1118) ,
  \2613(444)  = ~\2607(358) ,
  \981(1377)  = \940(1318)  & (\967(1204)  & (\930(1317)  & (\949(1369)  & \957(1370) ))),
  \271(181)  = \IN-271(181) ,
  \2470(456)  = ~\2468(373)  | ~\2461(285) ,
  \2018(404)  = ~\2012(313) ,
  \1934(980)  = \1912(959)  & \1994(267) ,
  \2099(249)  = ~\2096(218) ,
  \1025(1399)  = \487(403)  & \644(1391) ,
  \1213(585)  = ~\1470(562)  | ~\2099(249) ,
  \2370(1192)  = ~\2366(1132) ,
  \897(755)  = \889(670)  | \887(597) ,
  \2175(871)  = ~\2169(782) ,
  \1861(1049)  = \1842(1037)  & \2094(251) ,
  \999(895)  = ~\995(798) ,
  \164(607)  = \[104] ,
  \1085(1408)  = \1830(1108)  & (\1027(1407)  & \690(1393) ),
  \1742(530)  = \1728(406)  & \21(14) ,
  \2141(793)  = \1080(705) ,
  \219(302)  = \[85] ,
  \2705(339)  = ~\2699(248) ,
  \824(508)  = \795(294)  & (\784(378)  & \56(41) ),
  \2550(835)  = ~\2546(743) ,
  \1754(854)  = ~\1753(674)  | ~\1752(762) ,
  \335(299)  = \452(190) ,
  \967(1204)  = \1051(695)  & \1382(1116) ,
  \547(415)  = ~\546(322) ,
  \1449(467)  = \1430(336)  & (\1406(338)  & \136(107) ),
  \2034(633)  = \2012(313)  & \1464(560) ,
  \1307(492)  = \1296(374)  & (\1273(377)  & \89(68) ),
  \633(1142)  = \617(1077)  & (\575(1021)  & \584(1074) ),
  \1087(1275)  = ~\1093(1220) ,
  \1524(579)  = ~\1521(541) ,
  \456(709)  = \40(29)  & (\1387(594)  & \1389(610) ),
  \1164(1169)  = \708(1104)  & \1943(1097) ,
  \2766(808)  = ~\2762(716) ,
  \2371(1160)  = \1949(1090) ,
  \687(1357)  = ~\686(1329) ,
  \650(1380)  = ~\649(1346)  | ~\648(1366) ,
  \1118(1274)  = ~\2362(1194)  | ~\2355(1162) ,
  \1182(1343)  = ~\1181(1261)  | ~\1180(1313) ,
  \2639(605)  = \1704(557) ,
  \2551(372)  = \1344(286) ,
  \972(1347)  = \910(1301)  & (\924(1151)  & (\901(1303)  & \918(1305) )),
  \2565(455)  = ~\2559(370) ,
  \1317(459)  = \1284(293)  & \1273(377) ,
  \1475(331)  = ~\2433(242)  | ~\2430(224) ,
  \2541(902)  = ~\2535(825) ,
  \882(317)  = \868(198)  & \11(8) ,
  \2581(452)  = ~\2575(366) ,
  \1872(979)  = \1850(956)  & \1994(267) ,
  \2759(345)  = \2082(255) ,
  \819(509)  = \807(375)  & (\772(297)  & \55(40) ),
  \2775(341)  = \2094(251) ,
  \2524(576)  = ~\2522(539)  | ~\2515(553) ,
  \2310(1173)  = \534(1100) ,
  \922(1137)  = \499(1072)  & \1887(1086) ,
  \1689(381)  = \1655(243)  & (\1631(245)  & \117(92) ),
  \235(307)  = \[88] ,
  \1189(1348)  = \1128(1302)  & (\1142(1153)  & (\1119(1304)  & \1136(1306) )),
  \1568(1005)  = ~\1567(920) ,
  \202(139)  = \IN-202(139) ,
  \609(867)  = ~\2176(776)  | ~\2169(782) ,
  \1454(486)  = \1430(336)  & (\1394(246)  & \99(76) ),
  \177(116)  = \IN-177(116) ,
  \1323(496)  = \1296(374)  & (\1273(377)  & \85(64) ),
  \2390(1178)  = \714(1105) ,
  \2782(804)  = ~\2778(711) ,
  \2138(880)  = ~\2134(787) ,
  \1856(1051)  = \1842(1037)  & \2088(253) ,
  \1316(515)  = \1296(374)  & (\1261(296)  & \49(34) ),
  \1072(628)  = \1333(571) ,
  \2158(708)  = ~\2154(631) ,
  \1335(572)  = \1326(398)  | (\1325(505)  | (\1324(517)  | \1323(496) )),
  \244(158)  = \IN-244(158) ,
  \571(929)  = ~\570(890)  | ~\569(864) ,
  \2673(769)  = ~\2671(658)  | ~\2668(614) ,
  \239(153)  = \IN-239(153) ,
  \2205(1147)  = ~\2203(1081)  | ~\2200(1031) ,
  \2056(830)  = ~\2774(805)  | ~\2767(343) ,
  \823(518)  = \807(375)  & (\772(297)  & \43(30) ),
  \2318(1231)  = \528(1172) ,
  \1106(1201)  = \1035(618)  & \1624(1120) ,
  \2185(940)  = ~\2183(883)  | ~\2180(788) ,
  \2281(1212)  = ~\2275(1155) ,
  \1745(641)  = \1721(315)  & \1329(569) ,
  \208(145)  = \IN-208(145) ,
  \255(169)  = \IN-255(169) ,
  \218(311)  = \[84] ,
  \1762(764)  = ~\2646(675)  | ~\2639(605) ,
  \2225(1148)  = ~\2223(1082)  | ~\2220(1032) ,
  \2361(1219)  = ~\2355(1162) ,
  \552(460)  = \1256(401)  & \567(194) ,
  \613(1078)  = \589(1026) ,
  \1371(1056)  = \1361(1038)  & \2076(257) ,
  \199(136)  = \IN-199(136) ,
  \1794(430)  = ~\2698(344)  | ~\2691(252) ,
  \1643(337)  = ~\1631(245) ,
  \266(176)  = \IN-266(176) ,
  \605(1022)  = ~\601(930) ,
  \592(760)  = \562(672) ,
  \1227(681)  = \1470(562)  & \1213(585) ,
  \1885(1087)  = \1845(953)  & \1870(982) ,
  \1573(751)  = ~\2581(452)  | ~\2578(726) ,
  \1925(992)  = \1898(958)  & \1974(275) ,
  \988(1387)  = ~\969(1359)  | ~\976(1373) ,
  \1273(377)  = ~\1261(296) ,
  \2338(873)  = ~\2334(784) ,
  \1828(1048)  = ~\2733(961)  | ~\2730(546) ,
  \2750(809)  = ~\2746(717) ,
  \2535(825)  = ~\1539(732)  | ~\1542(731) ,
  \277(187)  = \IN-277(187) ,
  \1074(703)  = ~\1072(628) ,
  \2401(1227)  = ~\2395(1170) ,
  \1748(534)  = \1728(406)  & \6(5) ,
  \473(1420)  = \1247(1418)  | \471(1419) ,
  \1826(1299)  = ~\2725(1247)  | ~\2722(1047) ,
  \2586(722)  = \1743(642)  | \1742(530) ,
  \1584(993)  = ~\1583(916) ,
  \1560(1221)  = \894(533)  & (\1559(1109)  & \1556(1111) ),
  \2076(257)  = ~\2072(214) ,
  \323(923)  = \896(846) ,
  \369(289)  = \1083(199) ,
  \579(866)  = ~\2122(774)  | ~\2115(780) ,
  \282(922)  = \896(846) ,
  \1156(1297)  = ~\2401(1227)  | ~\2398(1177) ,
  \896(846)  = \886(757)  | \885(596) ,
  \807(375)  = ~\795(294) ,
  \1326(398)  = \1284(293)  & (\1261(296)  & \72(53) ),
  \1945(1096)  = \1893(410)  & \1930(986) ,
  \1117(1251)  = ~\2361(1219)  | ~\2358(1136) ,
  \1035(618)  = ~\846(565) ,
  \1864(1112)  = \1863(991)  | \1861(1049) ,
  \2027(525)  = \2007(405)  & \26(19) ,
  \1457(425)  = \1430(336)  & \1406(338) ,
  \826(489)  = \807(375)  & (\784(378)  & \92(71) ),
  \575(1021)  = ~\571(929) ,
  \2478(234)  = ~\2474(231) ,
  \1692(472)  = \1655(243)  & (\1643(337)  & \128(101) ),
  \2650(606)  = \1707(558) ,
  \690(1393)  = ~\688(1381) ,
  \642(1345)  = ~\2234(1263)  | ~\2227(1308) ,
  \947(1353)  = ~\2321(1320)  | ~\2318(1231) ,
  \2716(928)  = ~\2712(861) ,
  \1148(1323)  = ~\1147(1283)  | ~\1146(1298) ,
  \2654(677)  = ~\2650(606) ,
  \1801(1017)  = ~\1798(927) ,
  \2468(373)  = ~\2464(287) ,
  \2347(1185)  = \1624(1120) ,
  \1368(1058)  = \1361(1038)  & \2070(260) ,
  \525(1029)  = \769(878)  | \767(937) ,
  \1146(1298)  = ~\2393(1226)  | ~\2390(1178) ,
  \743(800)  = ~\456(709) ,
  \1594(837)  = ~\2622(811)  | ~\2615(356) ,
  \2403(1285)  = \1941(1228) ,
  \971(1336)  = \922(1137)  & (\901(1303)  & \910(1301) ),
  \1078(629)  = \1335(572) ,
  \1575(918)  = ~\1574(842)  | ~\1573(751) ,
  \2267(1158)  = \1891(1088) ,
  \303(698)  = \1060(626) ,
  \2062(968)  = ~\2061(906) ,
  \1194(1383)  = \1175(1372)  & (\1148(1323)  & (\1167(1371)  & (\1182(1343)  & \1158(1324) ))),
  \2040(834)  = ~\2742(807)  | ~\2735(352) ,
  \1389(610)  = ~\1464(560) ,
  \948(1319)  = ~\2322(1290)  | ~\2315(1281) ,
  \2059(736)  = ~\2781(429)  | ~\2778(711) ,
  \1555(1064)  = \1564(1008)  & (\1568(1005)  & (\1572(1002)  & (\1576(999)  & \1580(996) ))),
  \2503(445)  = ~\2501(357)  | ~\2498(272) ,
  \1256(401)  = ~\1254(308) ,
  \701(1103)  = \994(412)  & \699(1030) ,
  \492(1035)  = \742(951)  & \490(886) ,
  \588(936)  = ~\2130(875)  | ~\2123(697) ,
  \2697(342)  = ~\2691(252) ,
  \1553(1110)  = ~\1552(978)  | ~\1551(1062) ,
  \1509(552)  = ~\1508(451)  | ~\1507(453) ,
  \409(298)  = \452(190) ,
  \1310(394)  = \1284(293)  & (\1261(296)  & \76(57) ),
  \2043(741)  = ~\2749(437)  | ~\2746(717) ,
  \954(1289)  = \528(1172)  & \1879(1224) ,
  \1521(541)  = \1495(419) ,
  \2210(933)  = ~\2160(778)  | ~\2159(892) ,
  \881(408)  = \875(290)  & \11(8) ,
  \1158(1324)  = ~\1157(1284)  | ~\1156(1297) ,
  \2533(664)  = ~\2531(589)  | ~\2528(550) ,
  \183(122)  = \IN-183(122) ,
  \830(490)  = \807(375)  & (\784(378)  & \91(70) ),
  \2554(724)  = \1735(645)  | \1734(532) ,
  \2190(792)  = \1074(703) ,
  \250(164)  = \IN-250(164) ,
  \1394(246)  = \2104(220) ,
  \1250(604)  = \1704(557) ,
  \1188(1337)  = \1140(1139)  & (\1119(1304)  & \1128(1302) ),
  \2323(1282)  = \1877(1225) ,
  \1827(1238)  = ~\2726(1107)  | ~\2719(1190) ,
  \2726(1107)  = ~\2722(1047) ,
  \2570(723)  = \1739(647)  | \1738(531) ,
  \2715(904)  = ~\2709(827) ,
  \2224(1080)  = ~\2220(1032) ,
  \234(376)  = \[97] ,
  \2374(1140)  = \726(1073) ,
  \639(1126)  = \625(1076)  & (\596(853)  & \605(1022) ),
  \2114(771)  = ~\2110(685) ,
  \2103(247)  = ~\2100(219) ,
  \2024(636)  = \2001(314)  & \1698(563) ,
  \1818(1011)  = \1802(926)  & (\1758(924)  & \1767(925) ),
  \2738(714)  = \2026(639)  | \2025(522) ,
  \1591(914)  = ~\1590(838)  | ~\1589(746) ,
  \1378(1121)  = \1369(1004)  | \1368(1058) ,
  \1578(841)  = ~\2590(814)  | ~\2583(364) ,
  \2157(777)  = ~\2151(691) ,
  \1127(1271)  = ~\2370(1192)  | ~\2363(1159) ,
  \272(182)  = \IN-272(182) ,
  \1507(453)  = ~\2485(365)  | ~\2482(280) ,
  \898(756)  = \893(598)  | \891(669) ,
  \194(131)  = \IN-194(131) ,
  \2706(340)  = ~\2702(250) ,
  \1687(480)  = \1667(334)  & (\1631(245)  & \105(82) ),
  \725(1020)  = \1005(952)  & \723(863) ,
  \1173(1354)  = ~\2417(1328)  | ~\2414(1234) ,
  \321(848)  = \897(755) ,
  \1863(991)  = \1836(955)  & \1974(275) ,
  \1119(1304)  = ~\1118(1274)  | ~\1117(1251) ,
  \833(392)  = \795(294)  & (\772(297)  & \78(59) ),
  \2614(817)  = ~\2610(725) ,
  \490(886)  = \743(800)  & \1078(629) ,
  \1877(1225)  = \1831(409)  & \1859(1114) ,
  \1544(651)  = \1529(592)  & (\1500(538)  & \1509(552) ),
  \2123(697)  = ~\1057(624) ,
  \1261(296)  = \543(192) ,
  \2754(713)  = \2030(637)  | \2029(521) ,
  \708(1104)  = ~\707(1043) ,
  \203(140)  = \IN-203(140) ,
  \748(411)  = \655(319) ,
  \1406(338)  = ~\1394(246) ,
  \2168(772)  = ~\2164(686) ,
  \2709(827)  = ~\2674(734)  | ~\2673(769) ,
  \1500(538)  = ~\1499(324)  | ~\1498(417) ,
  \2514(439)  = ~\2512(355)  | ~\2505(266) ,
  \937(1163)  = \540(1101)  & \1883(1094) ,
  \2487(274)  = \1976(207) ,
  \980(1384)  = \940(1318)  & (\961(1288)  & (\930(1317)  & \949(1369) )),
  \2387(1168)  = \1945(1096) ,
  \1920(995)  = \1898(958)  & \1969(277) ,
  \1147(1283)  = ~\2394(1237)  | ~\2387(1168) ,
  \2663(767)  = ~\2661(680)  | ~\2658(611) ,
  \337(263)  = \2066(212) ,
  \2770(712)  = \2034(633)  | \2033(520) ,
  \2204(1079)  = ~\2200(1031) ,
  \2712(861)  = ~\2664(768)  | ~\2663(767) ,
  \649(1346)  = ~\2250(1264)  | ~\2243(1300) ,
  \1682(469)  = \1667(334)  & (\1643(337)  & \131(104) ),
  \968(1333)  = \901(1303)  & (\918(1305)  & (\927(1315)  & \910(1301) )),
  \155(967)  = \1243(828)  | \1096(905) ,
  \1455(477)  = \1418(244)  & (\1406(338)  & \123(96) ),
  \1495(419)  = ~\1494(328)  | ~\1493(327) ,
  \795(294)  = \651(195) ,
  \2757(435)  = ~\2751(347) ,
  \1784(436)  = ~\2689(346)  | ~\2686(258) ,
  \957(1370)  = ~\956(1321)  | ~\955(1351) ,
  \2615(356)  = \1989(269) ,
  \1786(548)  = ~\1785(434)  | ~\1784(436) ,
  \1180(1313)  = ~\2425(1240)  | ~\2422(783) ,
  \256(170)  = \IN-256(170) ,
  \236(303)  = \[89] ,
  \749(801)  = \456(709) ,
  \769(878)  = \749(801)  & \1060(626) ,
  \2773(431)  = ~\2767(343) ,
  \1016(938)  = \999(895)  & \1060(626) ,
  \1776(323)  = ~\2682(233)  | ~\2675(261) ,
  \2065(715)  = \2038(635)  | \2037(523) ,
  \2322(1290)  = ~\2318(1231) ,
  \732(1068)  = ~\731(1013) ,
  \1541(577)  = \1525(540)  & (\1481(543)  & \1490(542) ),
  \1380(1118)  = \1373(1000)  | \1371(1056) ,
  \2046(974)  = ~\2045(910) ,
  \978(1349)  = \946(1165)  & \930(1317) ,
  \1752(762)  = ~\2637(683)  | ~\2634(555) ,
  \2307(1166)  = \1881(1095) ,
  \1735(645)  = \1710(316)  & \841(573) ,
  \1452(386)  = \1418(244)  & (\1394(246)  & \112(87) ),
  \1476(332)  = ~\2434(241)  | ~\2427(223) ,
  \1113(1368)  = \1110(1211)  & (\1100(1341)  & \1112(1339) ),
  \229(1180)  = \[128] ,
  \2485(365)  = ~\2479(278) ,
  \504(1012)  = \742(951)  & \502(855) ,
  \2337(1239)  = ~\2331(1181) ,
  \2630(810)  = ~\2626(718) ,
  \259(414)  = \[93] ,
  \1057(624)  = \1327(568) ,
  \1157(1284)  = ~\2402(1236)  | ~\2395(1170) ,
  \2241(770)  = ~\2235(684) ,
  \1858(994)  = \1836(955)  & \1969(277) ,
  \1344(286)  = ~\1341(200) ,
  \2471(282)  = \1956(203) ,
  \487(403)  = ~\486(312) ,
  \887(597)  = \875(290)  & \846(565) ,
  \325(507)  = \558(400) ,
  \1107(1061)  = \1607(1040)  & \1999(265) ,
  \940(1318)  = ~\939(1280)  | ~\938(1291) ,
  \1738(531)  = \1716(407)  & \20(13) ,
  \551(544)  = ~\550(422) ,
  \2538(730)  = ~\2524(576)  | ~\2523(653) ,
  \930(1317)  = ~\929(1279)  | ~\928(1292) ,
  \1704(557)  = \1693(382)  | (\1692(472)  | (\1691(481)  | \1690(463) )),
  \1751(643)  = \1721(315)  & \1335(572) ,
  \1140(1139)  = \726(1073)  & \1949(1090) ,
  \1199(1395)  = \1198(1378)  | (\1197(1385)  | (\1196(1355)  | (\1195(1350)  | \1155(1167) ))),
  \1080(705)  = ~\1078(629) ,
  \2082(255)  = ~\2078(215) ,
  \2460(326)  = ~\2458(235)  | ~\2451(229) ,
  \2498(272)  = \1981(208) ,
  \963(1262)  = ~\2338(873)  | ~\2331(1181) ,
  \2741(438)  = ~\2735(352) ,
  \178(117)  = \IN-178(117) ,
  \2457(236)  = ~\2451(229) ,
  \1193(1374)  = ~\1190(1362) ,
  \2186(944)  = ~\2184(881)  | ~\2177(790) ,
  \245(159)  = \IN-245(159) ,
  \1562(845)  = ~\2558(816)  | ~\2551(372) ,
  \767(937)  = \753(896)  & \1060(626) ,
  \1319(495)  = \1296(374)  & (\1273(377)  & \86(65) ),
  \1597(744)  = ~\2629(440)  | ~\2626(718) ,
  \1825(821)  = ~\1824(650)  & ~\1823(728) ,
  \977(1382)  = \957(1370)  & (\930(1317)  & (\949(1369)  & (\964(1344)  & \940(1318) ))),
  \2297(1214)  = ~\2291(1157) ,
  \2001(314)  = \29(22) ,
  \176(803)  = \[109] ,
  \189(126)  = \IN-189(126) ,
  \2441(240)  = ~\2435(225) ,
  \153(671)  = \[108] ,
  \927(1315)  = ~\926(1269)  | ~\925(1265) ,
  \2033(520)  = \2018(404)  & \34(25) ,
  \516(616)  = \838(564) ,
  \674(1200)  = \1035(618)  & \1378(1121) ,
  \894(533)  = \882(317)  | \881(408) ,
  \1321(504)  = \1284(293)  & (\1273(377)  & \61(44) ),
  \836(501)  = \795(294)  & (\784(378)  & \64(47) ),
  \2053(908)  = ~\2052(831)  | ~\2051(738) ,
  \608(932)  = ~\2175(871)  | ~\2172(690) ,
  \2671(658)  = ~\2665(582) ,
  \267(177)  = \IN-267(177) ,
  \1607(1040)  = ~\1601(960) ,
  \2298(1208)  = ~\2294(1152) ,
  \2377(1217)  = ~\2371(1160) ,
  \1142(1153)  = \1947(1091)  & \720(1084) ,
  \1836(955)  = \475(897) ,
  \569(864)  = ~\2113(795)  | ~\2110(685) ,
  \820(498)  = \795(294)  & (\784(378)  & \67(50) ),
  \1921(1115)  = \1920(995)  | \1918(1052) ,
  \1096(905)  = \1243(828)  & \1228(735) ,
  \1930(986)  = \1898(958)  & \1984(271) ,
  \2482(280)  = \1961(204) ,
  \1460(335)  = \1418(244)  & \1394(246) ,
  \329(1414)  = \1208(1412) ,
  \1554(1063)  = \1584(993)  & (\1588(990)  & (\1592(987)  & (\1596(984)  & \1600(981) ))),
  \209(146)  = \IN-209(146) ,
  \1100(1341)  = ~\1099(1259)  | ~\1098(1311) ,
  \1041(620)  = \854(566) ,
  \144(601)  = \860(197)  & \838(564) ,
  \278(188)  = \IN-278(188) ,
  \681(1340)  = ~\684(1258)  | ~\683(1310) ,
  \1614(1059)  = \1607(1040)  & \2070(260) ,
  \213(150)  = \IN-213(150) ,
  \696(1175)  = ~\695(1102) ,
  \2226(1150)  = ~\2224(1080)  | ~\2217(1034) ,
  \2257(1241)  = ~\2251(1183) ,
  \1581(748)  = ~\2597(448)  | ~\2594(721) ,
  \1559(1109)  = \1558(1053)  & \1557(1093) ,
  \738(1071)  = ~\737(1015) ,
  \2668(614)  = \1470(562) ,
  \2203(1081)  = ~\2197(1033) ,
  \188(761)  = \[110] ,
  \546(322)  = \3(2)  & \1(0) ,
  \2223(1082)  = ~\2217(1034) ,
  \2012(313)  = \29(22) ,
  \970(1332)  = \915(1129)  & \901(1303) ,
  \231(1422)  = \[137] ,
  \220(306)  = \[86] ,
  \1569(752)  = ~\2573(454)  | ~\2570(723) ,
  \1955(320)  = \661(196)  & \7(6) ,
  \496(862)  = \743(800)  & \1698(563) ,
  \511(1070)  = ~\510(1014) ,
  \578(931)  = ~\2121(869)  | ~\2118(688) ,
  \901(1303)  = ~\900(1270)  | ~\899(1250) ,
  \160(609)  = \[102] ,
  \297(849)  = \898(756) ,
  \1445(466)  = \1430(336)  & (\1406(338)  & \137(108) ),
  \1814(1069)  = \1801(1017)  & (\1763(857)  & \1758(924) ),
  \2522(539)  = ~\2518(418) ,
  \1868(985)  = \1836(955)  & \1984(271) ,
  \1450(485)  = \1430(336)  & (\1394(246)  & \100(77) ),
  \2115(780)  = \1043(693) ,
  \1936(976)  = \1912(959)  & \1999(265) ,
  \1481(543)  = ~\1477(421) ,
  \2172(690)  = \1035(618) ,
  \2504(443)  = ~\2502(359)  | ~\2495(270) ,
  \2030(637)  = \2001(314)  & \1707(558) ,
  \2088(253)  = ~\2084(216) ,
  \1187(1334)  = \1133(1131)  & \1119(1304) ,
  \835(512)  = \807(375)  & (\772(297)  & \52(37) ),
  \1254(308)  = \69(52)  & (\108(85)  & (\57(42)  & \120(95) )),
  \2523(653)  = ~\2521(595)  | ~\2518(418) ,
  \1128(1302)  = ~\1127(1271)  | ~\1126(1249) ,
  \1228(735)  = \1227(681)  | \1225(660) ,
  \1504(575)  = ~\1500(538) ,
  \946(1165)  = \534(1100)  & \1881(1095) ,
  \1552(978)  = ~\2550(835)  | ~\2543(900) ,
  \1685(388)  = \1655(243)  & (\1631(245)  & \107(84) ),
  \1458(426)  = \1430(336)  & \1394(246) ,
  \1688(471)  = \1655(243)  & (\1643(337)  & \129(102) ),
  \240(154)  = \IN-240(154) ,
  \1234(657)  = \1473(545)  & \1218(583) ,
  \621(1075)  = \610(1024) ,
  \2515(553)  = ~\2470(456)  | ~\2469(458) ,
  \2698(344)  = ~\2694(254) ,
  \2534(663)  = ~\2532(590)  | ~\2525(549) ,
  \1744(529)  = \1728(406)  & \22(15) ,
  \184(123)  = \IN-184(123) ,
  \1296(374)  = ~\1284(293) ,
  \251(165)  = \IN-251(165) ,
  \2702(250)  = \2096(218) ,
  \2169(782)  = \1043(693) ,
  \1018(879)  = \995(798)  & \1060(626) ,
  \540(1101)  = ~\539(1042) ,
  \2200(1031)  = ~\2140(943)  | ~\2139(939) ,
  \195(132)  = \IN-195(132) ,
  \2306(1233)  = ~\2302(1174) ,
  \2220(1032)  = ~\2186(944)  | ~\2185(940) ,
  \1741(646)  = \1710(316)  & \857(567) ,
  \647(1307)  = ~\646(1254)  | ~\645(1197) ,
  \262(172)  = \IN-262(172) ,
  \2131(789)  = \1068(701) ,
  \2058(969)  = ~\2057(907) ,
  \2326(1230)  = \522(1171) ,
  \[100]  = ~\558(400) ,
  \1312(514)  = \1296(374)  & (\1261(296)  & \50(35) ),
  \918(1305)  = ~\917(1268)  | ~\916(1252) ,
  \2149(947)  = ~\2147(888)  | ~\2144(791) ,
  \628(1144)  = ~\625(1076) ,
  \1098(1311)  = ~\2345(1242)  | ~\2342(779) ,
  \[102]  = ~\1464(560) ,
  \2052(831)  = ~\2766(808)  | ~\2759(345) ,
  \1508(451)  = ~\2486(367)  | ~\2479(278) ,
  \2126(785)  = \1051(695) ,
  \2521(595)  = ~\2515(553) ,
  \[103]  = ~\1467(561) ,
  \1201(1398)  = \1200(1390)  | \1199(1395) ,
  \976(1373)  = ~\973(1361) ,
  \2531(589)  = ~\2525(549) ,
  \273(183)  = \IN-273(183) ,
  \1204(1405)  = ~\1201(1398) ,
  \[104]  = ~\1461(559) ,
  \693(1028)  = \1014(877)  | \1012(935) ,
  \1331(570)  = \1318(396)  | (\1317(459)  | (\1316(515)  | \1315(494) )),
  \596(853)  = ~\592(760) ,
  \[105]  = ~\1329(569) ,
  \2575(366)  = \1964(279) ,
  \1104(1203)  = \1043(693)  & \1626(1119) ,
  \2461(285)  = \1348(201) ,
  \[106]  = ~\1327(568) ,
  \2558(816)  = ~\2554(724) ,
  \631(1255)  = ~\630(1141)  & ~\629(1199) ,
  \1580(996)  = ~\1579(917) ,
  \[107]  = ~\857(567) ,
  \907(1133)  = \511(1070)  & \1891(1088) ,
  \493(1083)  = ~\492(1035) ,
  \[108]  = \152(599)  | \865(291) ,
  \899(1250)  = ~\2273(1215)  | ~\2270(1134) ,
  \[109]  = ~\175(710) ,
  \2508(268)  = \1991(210) ,
  \204(141)  = \IN-204(141) ,
  \2230(1206)  = ~\2206(1149)  | ~\2205(1147) ,
  \891(669)  = \875(290)  & \1041(620) ,
  \1184(1205)  = \1051(695)  & \1628(1117) ,
  \217(423)  = \[98] ,
  \2193(889)  = ~\2187(794) ,
  \2406(1235)  = \702(1176) ,
  \1999(265)  = ~\1996(211) ,
  \1051(695)  = ~\1049(622) ,
  \2039(742)  = ~\2741(438)  | ~\2738(714) ,
  \893(598)  = \868(198)  & \1327(568) ,
  \928(1292)  = ~\2305(1222)  | ~\2302(1174) ,
  \2197(1033)  = ~\2150(949)  | ~\2149(947) ,
  \246(160)  = \IN-246(160) ,
  \1953(1092)  = \1907(954)  & \1938(973) ,
  \[110]  = ~\187(673) ,
  \713(1044)  = \994(412)  & \711(946) ,
  \148(851)  = \[122] ,
  \1943(1097)  = \1893(410)  & \1928(989) ,
  \829(391)  = \795(294)  & (\772(297)  & \79(60) ),
  \1539(732)  = ~\1538(580)  & ~\1537(654) ,
  \938(1291)  = ~\2313(1223)  | ~\2310(1173) ,
  \2118(688)  = \1035(618) ,
  \1790(588)  = ~\1786(548) ,
  \1587(915)  = ~\1586(839)  | ~\1585(747) ,
  \2532(590)  = ~\2528(550) ,
  \2036(632)  = \2012(313)  & \1467(561) ,
  \2664(768)  = ~\2662(679)  | ~\2655(613) ,
  \257(171)  = \IN-257(171) ,
  \685(1375)  = \682(1367)  | (\680(1363)  | \671(1202) ),
  \498(1019)  = \742(951)  & \496(862) ,
  \521(1098)  = \748(411)  & \519(1027) ,
  \635(1189)  = \624(1143)  & (\601(930)  & \596(853) ),
  \290(704)  = \1078(629) ,
  \1823(728)  = \1813(661)  & (\1790(588)  & \1777(537) ),
  \2458(235)  = ~\2454(230) ,
  \471(1419)  = \1247(1418)  & \1240(1417) ,
  \2591(362)  = \1974(275) ,
  \2217(1034)  = ~\2196(950)  | ~\2195(948) ,
  \411(264)  = \2066(212) ,
  \2543(900)  = ~\1545(822)  | ~\1548(823) ,
  \1115(1257)  = ~\2354(773)  | ~\2347(1185) ,
  \2213(852)  = ~\2207(759) ,
  \1448(385)  = \1418(244)  & (\1394(246)  & \113(88) ),
  \2395(1170)  = \1943(1097) ,
  \1493(327)  = ~\2449(238)  | ~\2446(228) ,
  \1322(397)  = \1284(293)  & (\1261(296)  & \73(54) ),
  \720(1084)  = ~\719(1036) ,
  \2574(815)  = ~\2570(723) ,
  \1819(1128)  = ~\1818(1011)  & ~\1817(1066) ,
  \984(1397)  = \983(1389)  | \982(1394) ,
  \280(850)  = \898(756) ,
  \1785(434)  = ~\2690(348)  | ~\2683(256) ,
  \1615(1003)  = \1601(960)  & \1351(284) ,
  \1257(893)  = \468(797) ,
  \884(1386)  = \868(198)  & \650(1380) ,
  \2233(1338)  = ~\2227(1308) ,
  \2350(687)  = \1035(618) ,
  \2023(526)  = \2007(405)  & \25(18) ,
  \2151(691)  = ~\852(619) ,
  \2590(814)  = ~\2586(722) ,
  \2658(611)  = \1464(560) ,
  \2683(256)  = \2078(215) ,
  \[122]  = \147(600)  | \146(758) ,
  \237(309)  = \[90] ,
  \2342(779)  = \1043(693) ,
  \2418(1293)  = ~\2414(1234) ,
  \173(389)  = \[95] ,
  \955(1351)  = ~\2329(1322)  | ~\2326(1230) ,
  \2722(1047)  = ~\2718(965)  | ~\2717(1018) ,
  \1772(860)  = ~\1771(766)  | ~\1770(765) ,
  \2542(824)  = ~\2538(730) ,
  \909(1267)  = ~\2282(1191)  | ~\2275(1155) ,
  \1590(838)  = ~\2614(817)  | ~\2607(358) ,
  \[125]  = ~\155(967)  | ~\154(964) ,
  \2411(1286)  = \1939(1229) ,
  \1571(919)  = ~\1570(843)  | ~\1569(752) ,
  \179(118)  = \IN-179(118) ,
  \2055(737)  = ~\2773(431)  | ~\2770(712) ,
  \2618(719)  = \1751(643)  | \1750(527) ,
  \1166(1325)  = ~\2410(1296)  | ~\2403(1285) ,
  \1062(699)  = ~\1060(626) ,
  \[127]  = ~\1830(1108) ,
  \[128]  = ~\1553(1110) ,
  \2486(367)  = ~\2482(280) ,
  \480(292)  = \661(196) ,
  \1284(293)  = \651(195) ,
  \2275(1155)  = \1889(1085) ,
  \1830(1108)  = ~\1829(966)  | ~\1828(1048) ,
  \1874(975)  = \1850(956)  & \1999(265) ,
  \1678(461)  = \1667(334)  & (\1643(337)  & \142(113) ),
  \1747(640)  = \1721(315)  & \1331(570) ,
  \620(1145)  = ~\617(1077) ,
  \1859(1114)  = \1858(994)  | \1856(1051) ,
  \1798(927)  = \1772(860) ,
  \1631(245)  = \2104(220) ,
  \1135(1272)  = ~\2378(1196)  | ~\2371(1160) ,
  \2631(615)  = \1698(563) ,
  \630(1141)  = \613(1078)  & (\571(929)  & \580(1023) ),
  \1006(799)  = ~\456(709) ,
  \2274(1193)  = ~\2270(1134) ,
  \677(1122)  = \676(1006)  | \675(1060) ,
  \956(1321)  = ~\2330(1287)  | ~\2323(1282) ,
  \[130]  = ~\1560(1221) ,
  \1683(487)  = \1667(334)  & (\1631(245)  & \95(74) ),
  \910(1301)  = ~\909(1267)  | ~\908(1248) ,
  \1813(661)  = ~\1810(586) ,
  \[131]  = \144(601)  | \143(1330) ,
  \2661(680)  = ~\2655(613) ,
  \2645(676)  = ~\2639(605) ,
  \1031(630)  = ~\841(573) ,
  \308(1425)  = \1089(1423) ,
  \268(178)  = \IN-268(178) ,
  \1499(324)  = ~\2478(234)  | ~\2471(282) ,
  \533(1041)  = \748(411)  & \531(941) ,
  \1694(464)  = \1667(334)  & (\1643(337)  & \139(110) ),
  \846(565)  = \829(391)  | (\828(499)  | (\827(510)  | \826(489) )),
  \221(305)  = \[87] ,
  \1464(560)  = \1448(385)  | (\1447(475)  | (\1446(484)  | \1445(466) )),
  \158(349)  = \[92] ,
  \2094(251)  = ~\2090(217) ,
  \2743(350)  = \2070(260) ,
  \279(189)  = \IN-279(189) ,
  \[137]  = ~\473(1420) ,
  \1775(416)  = ~\2681(351)  | ~\2678(232) ,
  \214(151)  = \IN-214(151) ,
  \1824(650)  = \1810(586)  & (\1781(574)  & \1790(588) ),
  \929(1279)  = ~\2306(1233)  | ~\2299(1164) ,
  \1574(842)  = ~\2582(818)  | ~\2575(366) ,
  \[139]  = ~\1089(1423) ,
  \784(378)  = ~\772(297) ,
  \2559(370)  = \1351(284) ,
  \2029(521)  = \2007(405)  & \33(24) ,
  \331(1401)  = \895(1396) ,
  \1994(267)  = ~\1991(210) ,
  \2049(909)  = ~\2048(832)  | ~\2047(740) ,
  \1111(1364)  = \1106(1201)  & \1100(1341) ,
  \753(896)  = ~\749(801) ,
  \2196(950)  = ~\2194(885)  | ~\2187(794) ,
  \939(1280)  = ~\2314(1232)  | ~\2307(1166) ,
  \875(290)  = ~\868(198) ,
  \2605(446)  = ~\2599(360) ,
  \2602(720)  = \1747(640)  | \1746(528) ,
  \1200(1390)  = \1116(1376)  & \1194(1383) ,
  \2589(450)  = ~\2583(364) ,
  \857(567)  = \837(393)  | (\836(501)  | (\835(512)  | \834(491) )),
  \1459(424)  = \1418(244)  & \1406(338) ,
  \1093(1220)  = \14(9)  & \1092(1106) ,
  \2442(239)  = ~\2438(226) ,
  \2183(883)  = ~\2177(790) ,
  \1810(586)  = \1795(547) ,
  \2425(1240)  = ~\2419(1182) ,
  \1540(655)  = \1528(578)  & (\1490(542)  & \1477(421) ),
  \1750(527)  = \1728(406)  & \24(17) ,
  \2180(788)  = \1062(699) ,
  \1012(935)  = \999(895)  & \1057(624) ,
  \2694(254)  = \2084(216) ,
  \1005(952)  = \1257(893) ,
  \645(1197)  = ~\2241(770)  | ~\2238(1124) ,
  \1451(476)  = \1418(244)  & (\1406(338)  & \124(97) ),
  \2355(1162)  = \1953(1092) ,
  \2243(1300)  = ~\637(1245)  | ~\640(1246) ,
  \2672(682)  = ~\2668(614) ,
  \1543(750)  = \1532(666)  & (\1509(552)  & \1504(575) ),
  \2386(1209)  = ~\2382(1154) ,
  \1577(749)  = ~\2589(450)  | ~\2586(722) ,
  \1777(537)  = ~\1776(323)  | ~\1775(416) ,
  \1923(1050)  = \1904(1039)  & \2094(251) ,
  \765(876)  = \749(801)  & \1057(624) ,
  \895(1396)  = \884(1386)  | \883(668) ,
  \1989(269)  = ~\1986(209) ,
  \258(321)  = \661(196)  & (\15(10)  & \2(1) ),
  \1628(1117)  = \1623(998)  | \1621(1055) ,
  \241(155)  = \IN-241(155) ,
  \2557(457)  = ~\2551(372) ,
  \2345(1242)  = ~\2339(1184) ,
  \717(887)  = \1006(799)  & \1078(629) ,
  \190(127)  = \IN-190(127) ,
  \174(115)  = \IN-174(115) ,
  \1239(1415)  = \991(1411)  & \1221(1413) ,
  \1831(409)  = \658(318) ,
  \305(702)  = \1072(628) ,
  \2621(442)  = ~\2615(356) ,
  \2042(977)  = ~\2041(911) ,
  \1134(1253)  = ~\2377(1217)  | ~\2374(1140) ,
  \185(124)  = \IN-185(124) ,
  \2511(353)  = ~\2505(266) ,
  \686(1329)  = ~\1827(1238)  | ~\1826(1299) ,
  \2647(608)  = \1461(559) ,
  \2346(868)  = ~\2342(779) ,
  \2139(939)  = ~\2137(882)  | ~\2134(787) ,
  \146(758)  = \865(291)  & \562(672) ,
  \263(173)  = \IN-263(173) ,
  \1548(823)  = ~\1547(652)  & ~\1546(729) ,
  \2026(639)  = \2001(314)  & \1701(556) ,
  \196(133)  = \IN-196(133) ,
  \2758(806)  = ~\2754(713) ,
  \1734(532)  = \1716(407)  & \19(12) ,
  \2194(885)  = ~\2190(792) ,
  \1351(284)  = ~\1348(201) ,
  \1446(484)  = \1430(336)  & (\1394(246)  & \101(78) ),
  \2410(1296)  = ~\2406(1235) ,
  \171(621)  = \[107] ,
  \658(318)  = \8(7) ,
  \1315(494)  = \1296(374)  & (\1273(377)  & \87(66) ),
  \210(147)  = \IN-210(147) ,
  \841(573)  = \825(399)  | (\824(508)  | (\823(518)  | \822(497) )),
  \[84]  = ~\44(31) ,
  \1145(1316)  = ~\1144(1273)  | ~\1143(1266) ,
  \1373(1000)  = \1355(957)  & \1959(281) ,
  \1593(745)  = ~\2621(442)  | ~\2618(719) ,
  \[85]  = ~\132(105) ,
  \2385(1218)  = ~\2379(1161) ,
  \1533(591)  = \1518(551) ,
  \[86]  = ~\82(63) ,
  \617(1077)  = \589(1026) ,
  \169(114)  = \IN-169(114) ,
  \1125(1135)  = \738(1071)  & \1953(1092) ,
  \[87]  = ~\96(75) ,
  \205(142)  = \IN-205(142) ,
  \252(166)  = \IN-252(166) ,
  \[88]  = ~\69(52) ,
  \227(1179)  = \[127] ,
  \274(184)  = \IN-274(184) ,
  \1486(420)  = ~\1485(330)  | ~\1484(329) ,
  \1251(310)  = \44(31)  & (\96(75)  & (\82(63)  & \132(105) )),
  \[89]  = ~\120(95) ,
  \2573(454)  = ~\2567(368) ,
  \832(500)  = \795(294)  & (\784(378)  & \65(48) ),
  \763(934)  = \753(896)  & \1057(624) ,
  \1949(1090)  = \1907(954)  & \1934(980) ,
  \726(1073)  = ~\725(1020) ,
  \1387(594)  = \1385(283)  & \1461(559) ,
  \1327(568)  = \1310(394)  | (\1309(502)  | (\1308(513)  | \1307(492) )),
  \187(673)  = \547(415)  & (\554(581)  & (\483(191)  & \480(292) )),
  \166(625)  = \[105] ,
  \1737(648)  = \1710(316)  & \846(565) ,
  \223(413)  = \[96] ,
  \719(1036)  = \1005(952)  & \717(887) ,
  \1516(449)  = ~\2493(361)  | ~\2490(276) ,
  \636(1125)  = \621(1075)  & (\592(760)  & \601(930) ),
  \2187(794)  = \1080(705) ,
  \1596(984)  = ~\1595(913) ,
  \2235(684)  = \516(616) ,
  \2246(1207)  = ~\2226(1150)  | ~\2225(1148) ,
  \247(161)  = \IN-247(161) ,
  \[90]  = ~\57(42) ,
  \2294(1152)  = \493(1083) ,
  \1198(1378)  = \1158(1324)  & (\1184(1205)  & (\1148(1323)  & (\1167(1371)  & \1175(1372) ))),
  \[91]  = ~\108(85) ,
  \1904(1039)  = ~\1898(958) ,
  \2681(351)  = ~\2675(261) ,
  \1375(1054)  = \1361(1038)  & \2082(255) ,
  \961(1288)  = \522(1171)  & \1877(1225) ,
  \[92]  = ~\157(259) ,
  \2767(343)  = \2088(253) ,
  \1667(334)  = ~\1655(243) ,
  \2409(1326)  = ~\2403(1285) ,
  \2774(805)  = ~\2770(712) ,
  \[93]  = ~\258(321) ,
  \1889(1085)  = \1845(953)  & \1874(975) ,
  \2265(1244)  = ~\2259(1186) ,
  \1308(513)  = \1296(374)  & (\1261(296)  & \51(36) ),
  \2250(1264)  = ~\2246(1207) ,
  \2107(706)  = \1031(630) ,
  \531(941)  = \753(896)  & \1066(627) ,
  \1697(383)  = \1655(243)  & (\1631(245)  & \115(90) ),
  \[95]  = \654(300)  & \94(73) ,
  \1441(465)  = \1430(336)  & (\1406(338)  & \138(109) ),
  \589(1026)  = ~\588(936)  | ~\587(874) ,
  \[96]  = ~\1955(320) ,
  \[97]  = ~\1955(320)  | ~\567(194) ,
  \2144(791)  = \1074(703) ,
  \527(1099)  = \748(411)  & \525(1029) ,
  \[98]  = ~\216(333) ,
  \644(1391)  = ~\643(1379) ,
  \2329(1322)  = ~\2323(1282) ,
  \2578(726)  = \1741(646)  | \1740(535) ,
  \238(304)  = \[91] ,
  \2048(832)  = ~\2758(806)  | ~\2751(347) ,
  \924(1151)  = \1885(1087)  & \493(1083) ,
  \2045(910)  = ~\2044(833)  | ~\2043(741) ,
  \499(1072)  = ~\498(1019) ,
  \1144(1273)  = ~\2386(1209)  | ~\2379(1161) ,
  \2358(1136)  = \738(1071) ,
  \2238(1124)  = ~\2216(1065)  | ~\2215(1009) ,
  \1576(999)  = ~\1575(918) ,
  \2249(1331)  = ~\2243(1300) ,
  \1494(328)  = ~\2450(237)  | ~\2443(227) ,
  \1815(1010)  = \1798(927)  & (\1754(854)  & \1763(857) ),
  \2305(1222)  = ~\2299(1164) ,
  \1564(1008)  = ~\1563(921) ,
  \475(897)  = \462(802) ,
  \991(1411)  = \990(1402)  | \989(1409) ,
  \1565(753)  = ~\2565(455)  | ~\2562(727) ,
  \519(1027)  = \765(876)  | \763(934) ,
  \1770(765)  = ~\2653(678)  | ~\2650(606) ,
  \1802(926)  = \1772(860) ,
  \1805(1016)  = ~\1802(926) ,
  \286(696)  = \1057(624) ,
  \831(511)  = \807(375)  & (\772(297)  & \53(38) ),
  \1185(1335)  = \1119(1304)  & (\1136(1306)  & (\1145(1316)  & \1128(1302) )),
  \2742(807)  = ~\2738(714) ,
  \1926(1113)  = \1925(992)  | \1923(1050) ,
  \2254(781)  = \1043(693) ,
  \1258(894)  = \468(797) ,
  \1221(1413)  = ~\991(1411)  | ~\1208(1412) ,
  \1253(402)  = ~\1251(310) ,
  \1684(478)  = \1655(243)  & (\1643(337)  & \119(94) ),
  \2751(347)  = \2076(257) ,
  \2330(1287)  = ~\2326(1230) ,
  \550(422)  = \1253(402)  & \2106(222) ,
  \1470(562)  = \1456(387)  | (\1455(477)  | (\1454(486)  | \1453(468) )),
  \1324(517)  = \1296(374)  & (\1261(296)  & \47(32) ),
  \1599(912)  = ~\1598(836)  | ~\1597(744) ,
  \654(300)  = \452(190) ,
  \2314(1232)  = ~\2310(1173) ,
  \2781(429)  = ~\2775(341) ,
  \395(1392)  = \688(1381) ,
  \2150(949)  = ~\2148(884)  | ~\2141(793) ,
  \1883(1094)  = \1831(409)  & \1868(985) ,
  \865(291)  = ~\860(197) ,
  \2594(721)  = \1745(641)  | \1744(529) ,
  \666(1342)  = ~\665(1260)  | ~\664(1312) ,
  \2597(448)  = ~\2591(362) ,
  \587(874)  = ~\2129(786)  | ~\2126(785) ,
  \1318(396)  = \1284(293)  & (\1261(296)  & \74(55) ),
  \143(1330)  = \865(291)  & \647(1307) ,
  \1821(649)  = \1806(587)  & (\1777(537)  & \1786(548) ),
  \2394(1237)  = ~\2390(1178) ,
  \818(488)  = \807(375)  & (\784(378)  & \93(72) ),
  \1190(1362)  = \1189(1348)  | (\1188(1337)  | (\1187(1334)  | \1125(1135) )),
  \2689(346)  = ~\2683(256) ,
  \2354(773)  = ~\2350(687) ,
  \1136(1306)  = ~\1135(1272)  | ~\1134(1253) ,
  \915(1129)  = \505(1067)  & \1889(1085) ;
endmodule

