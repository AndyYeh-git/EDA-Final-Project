// IWLS benchmark module "C6288.iscas" printed on Wed May 29 16:29:58 2002
module test5 (\1GAT(0) , \18GAT(1) , \35GAT(2) , \52GAT(3) , \69GAT(4) , \86GAT(5) , \103GAT(6) , \120GAT(7) , \137GAT(8) , \154GAT(9) , \171GAT(10) , \188GAT(11) , \205GAT(12) , \222GAT(13) , \239GAT(14) , \256GAT(15) , \273GAT(16) , \290GAT(17) , \307GAT(18) , \324GAT(19) , \341GAT(20) , \358GAT(21) , \375GAT(22) , \392GAT(23) , \409GAT(24) , \426GAT(25) , \443GAT(26) , \460GAT(27) , \477GAT(28) , \494GAT(29) , \511GAT(30) , \528GAT(31) , \545GAT(287) , \1581GAT(423) , \1901GAT(561) , \2223GAT(700) , \2548GAT(840) , \2877GAT(983) , \3211GAT(1128) , \3552GAT(1275) , \3895GAT(1423) , \4241GAT(1572) , \4591GAT(1722) , \4946GAT(1876) , \5308GAT(2031) , \5672GAT(2187) , \5971GAT(2309) , \6123GAT(2368) , \6150GAT(2378) , \6160GAT(2383) , \6170GAT(2388) , \6180GAT(2393) , \6190GAT(2398) , \6200GAT(2403) , \6210GAT(2408) , \6220GAT(2413) , \6230GAT(2418) , \6240GAT(2423) , \6250GAT(2428) , \6260GAT(2433) , \6270GAT(2438) , \6280GAT(2443) , \6287GAT(2444) , \6288GAT(2447) );
input
  \137GAT(8) ,
  \154GAT(9) ,
  \443GAT(26) ,
  \103GAT(6) ,
  \171GAT(10) ,
  \120GAT(7) ,
  \188GAT(11) ,
  \409GAT(24) ,
  \494GAT(29) ,
  \69GAT(4) ,
  \18GAT(1) ,
  \86GAT(5) ,
  \35GAT(2) ,
  \460GAT(27) ,
  \52GAT(3) ,
  \477GAT(28) ,
  \1GAT(0) ,
  \324GAT(19) ,
  \341GAT(20) ,
  \307GAT(18) ,
  \392GAT(23) ,
  \358GAT(21) ,
  \511GAT(30) ,
  \375GAT(22) ,
  \528GAT(31) ,
  \222GAT(13) ,
  \239GAT(14) ,
  \205GAT(12) ,
  \290GAT(17) ,
  \256GAT(15) ,
  \273GAT(16) ,
  \426GAT(25) ;
output
  \6200GAT(2403) ,
  \3211GAT(1128) ,
  \3552GAT(1275) ,
  \6150GAT(2378) ,
  \545GAT(287) ,
  \1581GAT(423) ,
  \6270GAT(2438) ,
  \5308GAT(2031) ,
  \6287GAT(2444) ,
  \2223GAT(700) ,
  \6240GAT(2423) ,
  \6250GAT(2428) ,
  \6190GAT(2398) ,
  \5971GAT(2309) ,
  \2877GAT(983) ,
  \4946GAT(1876) ,
  \6220GAT(2413) ,
  \4241GAT(1572) ,
  \6160GAT(2383) ,
  \2548GAT(840) ,
  \6180GAT(2393) ,
  \5672GAT(2187) ,
  \6280GAT(2443) ,
  \3895GAT(1423) ,
  \6210GAT(2408) ,
  \4591GAT(1722) ,
  \6230GAT(2418) ,
  \6260GAT(2433) ,
  \1901GAT(561) ,
  \6123GAT(2368) ,
  \6170GAT(2388) ,
  \6288GAT(2447) ;
wire
  \4248GAT(1567) ,
  \2326GAT(742) ,
  \2591GAT(829) ,
  \4126GAT(1512) ,
  \1870GAT(518) ,
  \2467GAT(767) ,
  \603GAT(267) ,
  \1714GAT(440) ,
  \4278GAT(1556) ,
  \6177GAT(2389) ,
  \2024GAT(583) ,
  \4805GAT(1780) ,
  \1567GAT(371) ,
  \4215GAT(1525) ,
  \1533GAT(390) ,
  \4925GAT(1828) ,
  \6030GAT(2313) ,
  \2209GAT(645) ,
  \5617GAT(2162) ,
  \3145GAT(1094) ,
  \939GAT(155) ,
  \5785GAT(2231) ,
  \5374GAT(2056) ,
  \3784GAT(1359) ,
  \5254GAT(1994) ,
  \1621GAT(409) ,
  \4491GAT(1657) ,
  \1311GAT(302) ,
  \5428GAT(2083) ,
  \1450GAT(361) ,
  \4963GAT(1867) ,
  \1382GAT(321) ,
  \3496GAT(1247) ,
  \4901GAT(1845) ,
  \2611GAT(854) ,
  \4360GAT(1619) ,
  \4880GAT(1854) ,
  \2595GAT(858) ,
  \5052GAT(1894) ,
  \1946GAT(546) ,
  \1917GAT(555) ,
  \1871GAT(516) ,
  \1672GAT(428) ,
  \639GAT(255) ,
  \3486GAT(1251) ,
  \762GAT(214) ,
  \3410GAT(1177) ,
  \3921GAT(1411) ,
  \960GAT(148) ,
  \2856GAT(931) ,
  \5266GAT(1990) ,
  \4320GAT(1582) ,
  \4208GAT(1528) ,
  \5606GAT(2156) ,
  \4350GAT(1573) ,
  \5420GAT(2036) ,
  \5770GAT(2197) ,
  \3333GAT(1160) ,
  \3577GAT(1264) ,
  \5684GAT(2183) ,
  \681GAT(241) ,
  \4185GAT(1546) ,
  \774GAT(210) ,
  \3850GAT(1379) ,
  \6251GAT(2427) ,
  \1347GAT(293) ,
  \2151GAT(682) ,
  \3461GAT(1201) ,
  \3565GAT(1269) ,
  \5642GAT(2146) ,
  \5818GAT(2232) ,
  \1002GAT(134) ,
  \2269GAT(716) ,
  \6241GAT(2422) ,
  \2946GAT(997) ,
  \6037GAT(2332) ,
  \3170GAT(1082) ,
  \2857GAT(938) ,
  \4520GAT(1648) ,
  \3646GAT(1285) ,
  \5044GAT(1885) ,
  \2983GAT(984) ,
  \2245GAT(692) ,
  \846GAT(186) ,
  \5809GAT(2224) ,
  \5416GAT(2038) ,
  \1705GAT(450) ,
  \5251GAT(2004) ,
  \4727GAT(1759) ,
  \4428GAT(1644) ,
  \5747GAT(2205) ,
  \5676GAT(2185) ,
  \3253GAT(1119) ,
  \3015GAT(1013) ,
  \4698GAT(1727) ,
  \3052GAT(1040) ,
  \2028GAT(579) ,
  \5726GAT(2169) ,
  \2200GAT(655) ,
  \5688GAT(2191) ,
  \4791GAT(1784) ,
  \5192GAT(1968) ,
  \2150GAT(683) ,
  \5297GAT(1996) ,
  \3832GAT(1399) ,
  \4650GAT(1746) ,
  \3019GAT(1006) ,
  \1945GAT(545) ,
  \5013GAT(1900) ,
  \1355GAT(291) ,
  \4676GAT(1740) ,
  \2184GAT(657) ,
  \5030GAT(1891) ,
  \5022GAT(1898) ,
  \4359GAT(1610) ,
  \3425GAT(1214) ,
  \2011GAT(600) ,
  \5345GAT(2016) ,
  \861GAT(181) ,
  \4772GAT(1790) ,
  \804GAT(200) ,
  \4013GAT(1458) ,
  \3374GAT(1191) ,
  \4498GAT(1654) ,
  \3380GAT(1188) ,
  \5882GAT(2276) ,
  \6049GAT(2329) ,
  \4546GAT(1692) ,
  \3161GAT(1100) ,
  \3186GAT(1086) ,
  \2199GAT(648) ,
  \2029GAT(582) ,
  \1507GAT(407) ,
  \4800GAT(1782) ,
  \3687GAT(1301) ,
  \4845GAT(1809) ,
  \3103GAT(1063) ,
  \2185GAT(664) ,
  \2954GAT(995) ,
  \2201GAT(653) ,
  \1795GAT(492) ,
  \3202GAT(1080) ,
  \3437GAT(1211) ,
  \5332GAT(2033) ,
  \4064GAT(1486) ,
  \3536GAT(1230) ,
  \5618GAT(2161) ,
  \2558GAT(836) ,
  \1568GAT(369) ,
  \4922GAT(1829) ,
  \6256GAT(2431) ,
  \5472GAT(2061) ,
  \3524GAT(1225) ,
  \2089GAT(639) ,
  \3087GAT(1067) ,
  \4332GAT(1579) ,
  \3324GAT(1176) ,
  \4082GAT(1480) ,
  \4273GAT(1558) ,
  \4780GAT(1797) ,
  \5241GAT(2008) ,
  \2266GAT(684) ,
  \5544GAT(2134) ,
  \3926GAT(1420) ,
  \3046GAT(1042) ,
  \4646GAT(1747) ,
  \2516GAT(792) ,
  \3076GAT(1032) ,
  \5519GAT(2091) ,
  \3499GAT(1232) ,
  \3857GAT(1389) ,
  \2380GAT(757) ,
  \4519GAT(1647) ,
  \1315GAT(301) ,
  \2265GAT(686) ,
  \1594GAT(418) ,
  \3458GAT(1202) ,
  \3764GAT(1364) ,
  \1506GAT(406) ,
  \5645GAT(2145) ,
  \2777GAT(917) ,
  \597GAT(269) ,
  \5287GAT(1983) ,
  \876GAT(176) ,
  \6205GAT(2405) ,
  \5554GAT(2126) ,
  \1628GAT(439) ,
  \5813GAT(2233) ,
  \5911GAT(2264) ,
  \4509GAT(1651) ,
  \6010GAT(2323) ,
  \2410GAT(746) ,
  \4018GAT(1465) ,
  \4329GAT(1580) ,
  \2204GAT(646) ,
  \3835GAT(1384) ,
  \4203GAT(1529) ,
  \3932GAT(1408) ,
  \5275GAT(1988) ,
  \4159GAT(1499) ,
  \2980GAT(985) ,
  \4005GAT(1463) ,
  \4306GAT(1591) ,
  \3905GAT(1417) ,
  \4612GAT(1713) ,
  \594GAT(270) ,
  \2599GAT(857) ,
  \2603GAT(856) ,
  \3132GAT(1053) ,
  \4180GAT(1548) ,
  \4587GAT(1682) ,
  \5993GAT(2301) ,
  \3026GAT(1003) ,
  \4715GAT(1772) ,
  \1466GAT(357) ,
  \4634GAT(1704) ,
  \3398GAT(1182) ,
  \3336GAT(1169) ,
  \5840GAT(2257) ,
  \5427GAT(2076) ,
  \2414GAT(782) ,
  \4167GAT(1496) ,
  \1343GAT(294) ,
  \5366GAT(2058) ,
  \1547GAT(383) ,
  \5249GAT(1995) ,
  \5984GAT(2311) ,
  \3865GAT(1376) ,
  \4462GAT(1668) ,
  \5076GAT(1925) ,
  \4575GAT(1673) ,
  \5954GAT(2283) ,
  \2996GAT(1027) ,
  \3001GAT(1012) ,
  \1624GAT(408) ,
  \2671GAT(865) ,
  \2125GAT(630) ,
  \5439GAT(2080) ,
  \3847GAT(1393) ,
  \2905GAT(971) ,
  \3883GAT(1370) ,
  \2942GAT(998) ,
  \2273GAT(715) ,
  \2264GAT(685) ,
  \5063GAT(1879) ,
  \2021GAT(590) ,
  \5637GAT(2148) ,
  \2672GAT(872) ,
  \1296GAT(36) ,
  \1206GAT(66) ,
  \1077GAT(109) ,
  \1388GAT(315) ,
  \4398GAT(1596) ,
  \6246GAT(2426) ,
  \4620GAT(1710) ,
  \2582GAT(827) ,
  \2338GAT(730) ,
  \4118GAT(1514) ,
  \2191GAT(659) ,
  \5586GAT(2116) ,
  \4601GAT(1717) ,
  \4026GAT(1452) ,
  \3755GAT(1324) ,
  \5879GAT(2238) ,
  \4730GAT(1758) ,
  \5738GAT(2207) ,
  \2914GAT(967) ,
  \6108GAT(2362) ,
  \4160GAT(1507) ,
  \1299GAT(35) ,
  \1209GAT(65) ,
  \4977GAT(1863) ,
  \4947GAT(1875) ,
  \5522GAT(2090) ,
  \624GAT(260) ,
  \5526GAT(2088) ,
  \6157GAT(2379) ,
  \2186GAT(662) ,
  \4896GAT(1847) ,
  \4435GAT(1632) ,
  \1546GAT(382) ,
  \2781GAT(916) ,
  \5115GAT(1903) ,
  \2492GAT(817) ,
  \2190GAT(661) ,
  \5501GAT(2097) ,
  \1290GAT(38) ,
  \1293GAT(37) ,
  \1203GAT(67) ,
  \1200GAT(68) ,
  \5378GAT(2050) ,
  \5782GAT(2192) ,
  \4079GAT(1481) ,
  \546GAT(286) ,
  \6073GAT(2341) ,
  \6147GAT(2374) ,
  \2511GAT(795) ,
  \930GAT(158) ,
  \4838GAT(1816) ,
  \1437GAT(335) ,
  \2950GAT(996) ,
  \4531GAT(1698) ,
  \2242GAT(693) ,
  \3480GAT(1254) ,
  \1389GAT(314) ,
  \2917GAT(974) ,
  \4886GAT(1851) ,
  \1756GAT(469) ,
  \1351GAT(292) ,
  \2383GAT(756) ,
  \2649GAT(845) ,
  \2724GAT(894) ,
  \2339GAT(735) ,
  \1434GAT(336) ,
  \1597GAT(417) ,
  \2085GAT(640) ,
  \4189GAT(1545) ,
  \3453GAT(1204) ,
  \768GAT(212) ,
  \4985GAT(1861) ,
  \5870GAT(2242) ,
  \5611GAT(2155) ,
  \1011GAT(131) ,
  \4683GAT(1732) ,
  \1791GAT(493) ,
  \4174GAT(1551) ,
  \5262GAT(1992) ,
  \3501GAT(1245) ,
  \630GAT(258) ,
  \4708GAT(1768) ,
  \561GAT(281) ,
  \1390GAT(313) ,
  \5856GAT(2246) ,
  \849GAT(185) ,
  \5147GAT(1939) ,
  \5288GAT(1984) ,
  \1963GAT(573) ,
  \2670GAT(874) ,
  \2673GAT(864) ,
  \4907GAT(1834) ,
  \5080GAT(1916) ,
  \6045GAT(2334) ,
  \627GAT(259) ,
  \1044GAT(120) ,
  \2350GAT(719) ,
  \2113GAT(633) ,
  \3571GAT(1266) ,
  \6221GAT(2412) ,
  \1281GAT(41) ,
  \1221GAT(61) ,
  \3583GAT(1261) ,
  \2475GAT(765) ,
  \2493GAT(815) ,
  \1319GAT(300) ,
  \5430GAT(2082) ,
  \2023GAT(588) ,
  \2816GAT(949) ,
  \2861GAT(930) ,
  \2648GAT(842) ,
  \2189GAT(654) ,
  \1284GAT(40) ,
  \1224GAT(60) ,
  \3349GAT(1161) ,
  \5255GAT(2003) ,
  \3309GAT(1134) ,
  \2336GAT(732) ,
  \4739GAT(1754) ,
  \3146GAT(1106) ,
  \4760GAT(1795) ,
  \2555GAT(837) ,
  \4875GAT(1813) ,
  \1391GAT(312) ,
  \2337GAT(737) ,
  \2908GAT(970) ,
  \1287GAT(39) ,
  \1272GAT(44) ,
  \1227GAT(59) ,
  \1212GAT(64) ,
  \5483GAT(2103) ,
  \5837GAT(2252) ,
  \5996GAT(2300) ,
  \3697GAT(1297) ,
  \717GAT(229) ,
  \6119GAT(2358) ,
  \2666GAT(878) ,
  \2418GAT(781) ,
  \5845GAT(2256) ,
  \5476GAT(2075) ,
  \969GAT(145) ,
  \6135GAT(2369) ,
  \5395GAT(2045) ,
  \4837GAT(1812) ,
  \3162GAT(1099) ,
  \2790GAT(914) ,
  \1392GAT(311) ,
  \1384GAT(319) ,
  \4641GAT(1703) ,
  \2474GAT(764) ,
  \2811GAT(952) ,
  \4070GAT(1483) ,
  \1278GAT(42) ,
  \1218GAT(62) ,
  \2070GAT(610) ,
  \2481GAT(813) ,
  \3516GAT(1237) ,
  \3417GAT(1216) ,
  \1047GAT(119) ,
  \2727GAT(899) ,
  \4287GAT(1552) ,
  \714GAT(230) ,
  \3330GAT(1173) ,
  \4633GAT(1706) ,
  \1275GAT(43) ,
  \1215GAT(63) ,
  \4275GAT(1557) ,
  \5452GAT(2066) ,
  \4393GAT(1598) ,
  \4245GAT(1568) ,
  \4363GAT(1607) ,
  \3397GAT(1190) ,
  \1741GAT(475) ,
  \4849GAT(1807) ,
  \4525GAT(1701) ,
  \2813GAT(961) ,
  \933GAT(157) ,
  \5704GAT(2175) ,
  \5259GAT(1993) ,
  \4205GAT(1538) ,
  \4385GAT(1601) ,
  \1266GAT(46) ,
  \1236GAT(56) ,
  \4038GAT(1447) ,
  \3107GAT(1062) ,
  \2483GAT(820) ,
  \2022GAT(585) ,
  \5051GAT(1884) ,
  \5566GAT(2121) ,
  \4224GAT(1523) ,
  \5245GAT(2007) ,
  \3239GAT(1116) ,
  \1393GAT(310) ,
  \1385GAT(318) ,
  \2791GAT(912) ,
  \6076GAT(2340) ,
  \2334GAT(734) ,
  \5537GAT(2085) ,
  \4139GAT(1509) ,
  \3485GAT(1252) ,
  \1269GAT(45) ,
  \1239GAT(55) ,
  \3495GAT(1248) ,
  \5788GAT(2236) ,
  \3959GAT(1440) ,
  \3140GAT(1097) ,
  \5148GAT(1937) ,
  \1074GAT(110) ,
  \1911GAT(557) ,
  \2335GAT(739) ,
  \5715GAT(2172) ,
  \4710GAT(1766) ,
  \633GAT(257) ,
  \2491GAT(807) ,
  \3914GAT(1414) ,
  \3064GAT(1037) ,
  \1263GAT(47) ,
  \1260GAT(48) ,
  \1233GAT(57) ,
  \1230GAT(58) ,
  \3886GAT(1369) ,
  \4688GAT(1731) ,
  \6165GAT(2385) ,
  \1709GAT(446) ,
  \5109GAT(1906) ,
  \3034GAT(1048) ,
  \1257GAT(49) ,
  \1242GAT(54) ,
  \2353GAT(723) ,
  \1508GAT(405) ,
  \5312GAT(2028) ,
  \4354GAT(1622) ,
  \1577GAT(365) ,
  \2667GAT(869) ,
  \2482GAT(821) ,
  \4440GAT(1631) ,
  \3206GAT(1071) ,
  \3568GAT(1267) ,
  \3360GAT(1150) ,
  \1443GAT(333) ,
  \5902GAT(2266) ,
  \2301GAT(708) ,
  \3659GAT(1276) ,
  \5283GAT(1985) ,
  \3467GAT(1198) ,
  \6120GAT(2356) ,
  \2812GAT(962) ,
  \4860GAT(1804) ,
  \4091GAT(1476) ,
  \1248GAT(52) ,
  \1386GAT(317) ,
  \5127GAT(1944) ,
  \5157GAT(1935) ,
  \5510GAT(2107) ,
  \3302GAT(1135) ,
  \2020GAT(587) ,
  \741GAT(221) ,
  \1339GAT(295) ,
  \3645GAT(1282) ,
  \966GAT(146) ,
  \3454GAT(1207) ,
  \1562GAT(374) ,
  \2463GAT(770) ,
  \5336GAT(2020) ,
  \1245GAT(53) ,
  \5849GAT(2249) ,
  \4607GAT(1714) ,
  \1759GAT(470) ,
  \2644GAT(846) ,
  \3466GAT(1200) ,
  \4769GAT(1791) ,
  \4792GAT(1785) ,
  \5197GAT(1966) ,
  \3010GAT(1015) ,
  \4014GAT(1467) ,
  \3746GAT(1326) ,
  \1008GAT(132) ,
  \3063GAT(1043) ,
  \4200GAT(1540) ,
  \555GAT(283) ,
  \1176GAT(76) ,
  \1440GAT(334) ,
  \3120GAT(1059) ,
  \1576GAT(364) ,
  \687GAT(239) ,
  \4152GAT(1500) ,
  \819GAT(195) ,
  \1582GAT(422) ,
  \1548GAT(381) ,
  \879GAT(175) ,
  \2721GAT(895) ,
  \3014GAT(1008) ,
  \3826GAT(1402) ,
  \5206GAT(1962) ,
  \4879GAT(1842) ,
  \3975GAT(1432) ,
  \4704GAT(1725) ,
  \4994GAT(1872) ,
  \1502GAT(348) ,
  \549GAT(285) ,
  \5923GAT(2259) ,
  \3156GAT(1102) ,
  \1708GAT(445) ,
  \765GAT(213) ,
  \6185GAT(2395) ,
  \1387GAT(316) ,
  \1179GAT(75) ,
  \4549GAT(1681) ,
  \2665GAT(871) ,
  \6226GAT(2416) ,
  \4067GAT(1484) ,
  \6171GAT(2387) ,
  \1874GAT(511) ,
  \2664GAT(880) ,
  \3967GAT(1438) ,
  \3793GAT(1357) ,
  \5505GAT(2095) ,
  \3005GAT(1010) ,
  \4545GAT(1693) ,
  \3542GAT(1219) ,
  \4427GAT(1635) ,
  \945GAT(153) ,
  \2340GAT(728) ,
  \3136GAT(1058) ,
  \1707GAT(448) ,
  \4236GAT(1518) ,
  \1563GAT(372) ,
  \1173GAT(77) ,
  \1170GAT(78) ,
  \4671GAT(1741) ,
  \4989GAT(1874) ,
  \3181GAT(1089) ,
  \5486GAT(2101) ,
  \5907GAT(2273) ,
  \3650GAT(1280) ,
  \2588GAT(824) ,
  \1182GAT(74) ,
  \5072GAT(1926) ,
  \2073GAT(608) ,
  \5928GAT(2290) ,
  \5890GAT(2271) ,
  \2869GAT(928) ,
  \4916GAT(1844) ,
  \2462GAT(769) ,
  \4781GAT(1788) ,
  \843GAT(187) ,
  \5498GAT(2098) ,
  \2343GAT(731) ,
  \1446GAT(362) ,
  \4341GAT(1575) ,
  \2669GAT(867) ,
  \3296GAT(1140) ,
  \5514GAT(2093) ,
  \1735GAT(477) ,
  \4294GAT(1594) ,
  \4965GAT(1866) ,
  \1676GAT(427) ,
  \1188GAT(72) ,
  \3321GAT(1129) ,
  \3519GAT(1226) ,
  \6275GAT(2440) ,
  \1474GAT(355) ,
  \2498GAT(812) ,
  \1975GAT(570) ,
  \4941GAT(1823) ,
  \1700GAT(453) ,
  \3996GAT(1425) ,
  \4439GAT(1630) ,
  \5792GAT(2235) ,
  \5966GAT(2278) ,
  \4842GAT(1810) ,
  \6133GAT(2370) ,
  \1612GAT(412) ,
  \2821GAT(946) ,
  \1185GAT(73) ,
  \3510GAT(1242) ,
  \4488GAT(1658) ,
  \3329GAT(1164) ,
  \[10] ,
  \1706GAT(447) ,
  \4933GAT(1826) ,
  \[11] ,
  \1875GAT(515) ,
  \792GAT(204) ,
  \4817GAT(1821) ,
  \[12] ,
  \2040GAT(621) ,
  \5268GAT(1989) ,
  \2528GAT(794) ,
  \[13] ,
  \1979GAT(569) ,
  \4008GAT(1470) ,
  \[14] ,
  \2239GAT(694) ,
  \4130GAT(1511) ,
  \2868GAT(927) ,
  \[15] ,
  \3489GAT(1235) ,
  \2526GAT(789) ,
  \[16] ,
  \1879GAT(508) ,
  \1578GAT(363) ,
  \[17] ,
  \4314GAT(1589) ,
  \5225GAT(1956) ,
  \3943GAT(1405) ,
  \[18] ,
  \1161GAT(81) ,
  \6081GAT(2339) ,
  \[19] ,
  \2496GAT(804) ,
  \1701GAT(454) ,
  \807GAT(199) ,
  \5924GAT(2260) ,
  \1164GAT(80) ,
  \2991GAT(1022) ,
  \4766GAT(1792) ,
  \2631GAT(849) ,
  \750GAT(218) ,
  \3756GAT(1333) ,
  \2827GAT(956) ,
  \5916GAT(2262) ,
  \684GAT(240) ,
  \3150GAT(1091) ,
  \1561GAT(373) ,
  \3908GAT(1416) ,
  \2007GAT(604) ,
  \1829GAT(538) ,
  \1763GAT(500) ,
  \[20] ,
  \5460GAT(2078) ,
  \[21] ,
  \2342GAT(726) ,
  \3632GAT(1288) ,
  \6068GAT(2343) ,
  \[22] ,
  \1167GAT(79) ,
  \1152GAT(84) ,
  \1821GAT(484) ,
  \[23] ,
  \2043GAT(620) ,
  \3667GAT(1320) ,
  \3874GAT(1372) ,
  \1335GAT(296) ,
  \1876GAT(513) ,
  \1397GAT(306) ,
  \[24] ,
  \[25] ,
  \[26] ,
  \1702GAT(451) ,
  \[27] ,
  \5989GAT(2310) ,
  \2902GAT(973) ,
  \2668GAT(876) ,
  \5434GAT(2081) ,
  \[28] ,
  \2305GAT(707) ,
  \1820GAT(486) ,
  \[29] ,
  \2789GAT(913) ,
  \2006GAT(601) ,
  \1158GAT(82) ,
  \2181GAT(665) ,
  \4395GAT(1597) ,
  \2341GAT(733) ,
  \5399GAT(2043) ,
  \4377GAT(1603) ,
  \2488GAT(818) ,
  \1155GAT(83) ,
  \1704GAT(449) ,
  \5594GAT(2113) ,
  \6217GAT(2409) ,
  \3718GAT(1337) ,
  \[30] ,
  \948GAT(152) ,
  \3166GAT(1098) ,
  \2966GAT(989) ,
  \[31] ,
  \3305GAT(1138) ,
  \4365GAT(1606) ,
  \2180GAT(667) ,
  \4716GAT(1762) ,
  \4825GAT(1819) ,
  \1396GAT(307) ,
  \3592GAT(1259) ,
  \4572GAT(1674) ,
  \5560GAT(2124) ,
  \840GAT(188) ,
  \3199GAT(1072) ,
  \972GAT(144) ,
  \2395GAT(750) ,
  \2828GAT(954) ,
  \1738GAT(476) ,
  \5575GAT(2119) ,
  \5069GAT(1919) ,
  \1926GAT(552) ,
  \3079GAT(1069) ,
  \6089GAT(2353) ,
  \3734GAT(1331) ,
  \5607GAT(2166) ,
  \6031GAT(2314) ,
  \1703GAT(452) ,
  \2005GAT(605) ,
  \5193GAT(1973) ,
  \4394GAT(1609) ,
  \816GAT(196) ,
  \4432GAT(1633) ,
  \4668GAT(1736) ,
  \4034GAT(1449) ,
  \1660GAT(431) ,
  \5085GAT(1914) ,
  \1395GAT(308) ,
  \3675GAT(1316) ,
  \4754GAT(1750) ,
  \1197GAT(69) ,
  \1005GAT(133) ,
  \3804GAT(1349) ,
  \4420GAT(1636) ,
  \672GAT(244) ,
  \4450GAT(1627) ,
  \4921GAT(1843) ,
  \3603GAT(1256) ,
  \4216GAT(1526) ,
  \3955GAT(1441) ,
  \1880GAT(512) ,
  \558GAT(282) ,
  \5552GAT(2127) ,
  \5446GAT(2069) ,
  \5797GAT(2234) ,
  \4866GAT(1802) ,
  \2359GAT(717) ,
  \2587GAT(826) ,
  \6237GAT(2419) ,
  \2260GAT(687) ,
  \1462GAT(358) ,
  \3809GAT(1356) ,
  \3608GAT(1294) ,
  \1101GAT(101) ,
  \5354GAT(2014) ,
  \5267GAT(1991) ,
  \1826GAT(543) ,
  \5764GAT(2209) ,
  \3506GAT(1243) ,
  \4900GAT(1846) ,
  \621GAT(261) ,
  \1543GAT(384) ,
  \1478GAT(354) ,
  \3212GAT(1127) ,
  \2426GAT(779) ,
  \2358GAT(721) ,
  \873GAT(177) ,
  \1881GAT(510) ,
  \753GAT(217) ,
  \1753GAT(471) ,
  \4913GAT(1831) ,
  \2004GAT(603) ,
  \6046GAT(2330) ,
  \4598GAT(1719) ,
  \1394GAT(309) ,
  \1588GAT(420) ,
  \1401GAT(347) ,
  \3124GAT(1055) ,
  \2753GAT(923) ,
  \4358GAT(1620) ,
  \5021GAT(1893) ,
  \1542GAT(386) ,
  \2864GAT(929) ,
  \5919GAT(2261) ,
  \2277GAT(714) ,
  \5685GAT(2181) ,
  \5808GAT(2223) ,
  \2513GAT(803) ,
  \1017GAT(129) ,
  \6061GAT(2344) ,
  \5895GAT(2269) ,
  \4012GAT(1468) ,
  \4161GAT(1498) ,
  \591GAT(271) ,
  \5250GAT(2005) ,
  \1083GAT(107) ,
  \3637GAT(1287) ,
  \2257GAT(688) ,
  \1815GAT(487) ,
  \6056GAT(2326) ,
  \1191GAT(71) ,
  \5727GAT(2167) ,
  \5035GAT(1889) ,
  \702GAT(234) ,
  \4529GAT(1686) ,
  \1825GAT(544) ,
  \810GAT(198) ,
  \1194GAT(70) ,
  \5480GAT(2105) ,
  \4748GAT(1752) ,
  \870GAT(178) ,
  \1014GAT(130) ,
  \2502GAT(811) ,
  \5047GAT(1895) ,
  \5353GAT(2030) ,
  \2718GAT(896) ,
  \3676GAT(1304) ,
  \5608GAT(2165) ,
  \2586GAT(825) ,
  \3248GAT(1121) ,
  \3668GAT(1309) ,
  \2512GAT(805) ,
  \1331GAT(297) ,
  \795GAT(203) ,
  \4787GAT(1786) ,
  \2101GAT(636) ,
  \2236GAT(695) ,
  \6151GAT(2377) ,
  \1929GAT(551) ,
  \3515GAT(1239) ,
  \6267GAT(2434) ,
  \5344GAT(2018) ,
  \3841GAT(1396) ,
  \1750GAT(472) ,
  \1824GAT(541) ,
  \6141GAT(2373) ,
  \5734GAT(2213) ,
  \5709GAT(2189) ,
  \2785GAT(915) ,
  \1618GAT(410) ,
  \2913GAT(969) ,
  \2309GAT(706) ,
  \5861GAT(2255) ,
  \2398GAT(754) ,
  \4526GAT(1700) ,
  \1541GAT(385) ,
  \4049GAT(1444) ,
  \3091GAT(1066) ,
  \4677GAT(1734) ,
  \4298GAT(1593) ,
  \4122GAT(1513) ,
  \6018GAT(2318) ,
  \4508GAT(1660) ,
  \5240GAT(2009) ,
  \4318GAT(1583) ,
  \4110GAT(1516) ,
  \6255GAT(2430) ,
  \5426GAT(2084) ,
  \3190GAT(1076) ,
  \5471GAT(2060) ,
  \3527GAT(1224) ,
  \5829GAT(2216) ,
  \3917GAT(1413) ,
  \1116GAT(96) ,
  \2281GAT(713) ,
  \2503GAT(809) ,
  \2061GAT(614) ,
  \3037GAT(1047) ,
  \2117GAT(632) ,
  \3185GAT(1077) ,
  \3075GAT(1034) ,
  \5930GAT(2295) ,
  \6101GAT(2348) ,
  \2527GAT(796) ,
  \3067GAT(1036) ,
  \2230GAT(697) ,
  \2912GAT(968) ,
  \2497GAT(814) ,
  \2349GAT(725) ,
  \1571GAT(367) ,
  \4211GAT(1527) ,
  \906GAT(166) ,
  \1119GAT(95) ,
  \2573GAT(831) ,
  \2174GAT(663) ,
  \5759GAT(2200) ,
  \3000GAT(1023) ,
  \4863GAT(1803) ,
  \3620GAT(1291) ,
  \2470GAT(766) ,
  \5331GAT(2022) ,
  \1518GAT(399) ,
  \4621GAT(1723) ,
  \4812GAT(1777) ,
  \1113GAT(97) ,
  \1110GAT(98) ,
  \1585GAT(421) ,
  \2009GAT(602) ,
  \4859GAT(1814) ,
  \2749GAT(924) ,
  \3872GAT(1373) ,
  \5221GAT(1958) ,
  \4405GAT(1643) ,
  \1122GAT(94) ,
  \5878GAT(2240) ,
  \3227GAT(1122) ,
  \2794GAT(911) ,
  \4950GAT(1873) ,
  \3325GAT(1168) ,
  \6166GAT(2386) ,
  \5990GAT(2302) ,
  \1020GAT(128) ,
  \1080GAT(108) ,
  \2254GAT(689) ,
  \3215GAT(1126) ,
  \915GAT(163) ,
  \2348GAT(720) ,
  \3541GAT(1228) ,
  \3476GAT(1196) ,
  \5749GAT(2204) ,
  \3131GAT(1052) ,
  \5464GAT(2063) ,
  \4487GAT(1662) ,
  \5194GAT(1967) ,
  \5136GAT(1942) ,
  \1128GAT(92) ,
  \5065GAT(1921) ,
  \3257GAT(1110) ,
  \2049GAT(618) ,
  \5280GAT(1986) ,
  \6245GAT(2425) ,
  \1787GAT(494) ,
  \5531GAT(2104) ,
  \4696GAT(1728) ,
  \5124GAT(1946) ,
  \4613GAT(1711) ,
  \4998GAT(1856) ,
  \813GAT(197) ,
  \1399GAT(304) ,
  \5587GAT(2114) ,
  \4871GAT(1801) ,
  \4544GAT(1683) ,
  \1125GAT(93) ,
  \2176GAT(668) ,
  \3556GAT(1273) ,
  \4709GAT(1775) ,
  \2968GAT(988) ,
  \2008GAT(599) ,
  \5343GAT(2017) ,
  \4017GAT(1454) ,
  \5670GAT(2136) ,
  \615GAT(263) ,
  \6023GAT(2316) ,
  \2570GAT(832) ,
  \5886GAT(2275) ,
  \2517GAT(802) ,
  \909GAT(165) ,
  \2486GAT(810) ,
  \2870GAT(926) ,
  \1023GAT(127) ,
  \6064GAT(2346) ,
  \1831GAT(540) ,
  \3836GAT(1398) ,
  \1732GAT(478) ,
  \5693GAT(2190) ,
  \2175GAT(670) ,
  \1131GAT(91) ,
  \5867GAT(2243) ,
  \5081GAT(1924) ,
  \1640GAT(436) ,
  \5438GAT(2072) ,
  \1104GAT(100) ,
  \1573GAT(366) ,
  \4829GAT(1818) ,
  \1134GAT(90) ,
  \5324GAT(2023) ,
  \6070GAT(2342) ,
  \1398GAT(305) ,
  \2487GAT(819) ,
  \3337GAT(1158) ,
  \5612GAT(2164) ,
  \2501GAT(801) ,
  \6186GAT(2396) ,
  \6011GAT(2319) ,
  \3681GAT(1312) ,
  \4928GAT(1827) ,
  \2521GAT(790) ,
  \6128GAT(2365) ,
  \5348GAT(2032) ,
  \4099GAT(1485) ,
  \2967GAT(992) ,
  \3673GAT(1317) ,
  \3851GAT(1392) ,
  \4885GAT(1852) ,
  \5947GAT(2284) ,
  \4895GAT(1848) ,
  \1092GAT(104) ,
  \1819GAT(485) ,
  \2873GAT(932) ,
  \2663GAT(873) ,
  \5721GAT(2170) ,
  \2995GAT(1018) ,
  \552GAT(284) ,
  \2662GAT(882) ,
  \3815GAT(1346) ,
  \4530GAT(1699) ,
  \5713GAT(2173) ,
  \6085GAT(2355) ,
  \2522GAT(799) ,
  \4040GAT(1446) ,
  \5188GAT(1974) ,
  \2357GAT(718) ,
  \5218GAT(1959) ,
  \1668GAT(429) ,
  \1086GAT(106) ,
  \2179GAT(660) ,
  \5304GAT(1978) ,
  \1572GAT(368) ,
  \2076GAT(611) ,
  \2639GAT(844) ,
  \2233GAT(696) ,
  \3509GAT(1229) ,
  \4143GAT(1504) ,
  \2703GAT(903) ,
  \6197GAT(2399) ,
  \3805GAT(1350) ,
  \4680GAT(1733) ,
  \4389GAT(1611) ,
  \4984GAT(1860) ,
  \4043GAT(1457) ,
  \1830GAT(542) ,
  \2715GAT(898) ,
  \1050GAT(118) ,
  \1400GAT(303) ,
  \5494GAT(2108) ,
  \2222GAT(642) ,
  \2345GAT(729) ,
  \5234GAT(1954) ,
  \6082GAT(2337) ,
  \4175GAT(1550) ,
  \5289GAT(1982) ,
  \5935GAT(2293) ,
  \1694GAT(459) ,
  \2536GAT(787) ,
  \4264GAT(1560) ,
  \5873GAT(2241) ,
  \3604GAT(1295) ,
  \3165GAT(1083) ,
  \3582GAT(1263) ,
  \6196GAT(2401) ,
  \5101GAT(1909) ,
  \798GAT(202) ,
  \3147GAT(1105) ,
  \1146GAT(86) ,
  \2797GAT(910) ,
  \3986GAT(1429) ,
  \2507GAT(808) ,
  \3944GAT(1403) ,
  \2221GAT(641) ,
  \1615GAT(411) ,
  \2523GAT(797) ,
  \1695GAT(460) ,
  \759GAT(215) ,
  \3500GAT(1246) ,
  \4302GAT(1592) ,
  \6014GAT(2322) ,
  \3338GAT(1167) ,
  \885GAT(173) ,
  \3408GAT(1178) ,
  \3591GAT(1268) ,
  \1149GAT(85) ,
  \4178GAT(1536) ,
  \744GAT(220) ,
  \5804GAT(2225) ,
  \5844GAT(2251) ,
  \663GAT(247) ,
  \5639GAT(2147) ,
  \2745GAT(925) ,
  \1143GAT(87) ,
  \1140GAT(88) ,
  \2661GAT(875) ,
  \3559GAT(1272) ,
  \2660GAT(884) ,
  \6026GAT(2315) ,
  \3521GAT(1234) ,
  \1137GAT(89) ,
  \5740GAT(2206) ,
  \1470GAT(356) ,
  \2033GAT(580) ,
  \6281GAT(2442) ,
  \4571GAT(1687) ,
  \2365GAT(762) ,
  \4711GAT(1774) ,
  \5401GAT(2042) ,
  \5009GAT(1901) ,
  \4622GAT(1709) ,
  \1886GAT(507) ,
  \4225GAT(1533) ,
  \5213GAT(1961) ,
  \2826GAT(943) ,
  \3177GAT(1090) ,
  \3095GAT(1065) ,
  \1783GAT(495) ,
  \2344GAT(724) ,
  \1971GAT(571) ,
  \897GAT(169) ,
  \2822GAT(958) ,
  \5599GAT(2111) ,
  \5817GAT(2221) ,
  \942GAT(154) ,
  \5323GAT(2025) ,
  \1851GAT(528) ,
  \2962GAT(993) ,
  \5650GAT(2144) ,
  \2224GAT(699) ,
  \4055GAT(1490) ,
  \2347GAT(727) ,
  \4061GAT(1488) ,
  \5451GAT(2068) ,
  \4973GAT(1877) ,
  \4595GAT(1720) ,
  \1696GAT(457) ,
  \4335GAT(1578) ,
  \3401GAT(1181) ,
  \4073GAT(1493) ,
  \6032GAT(2312) ,
  \5858GAT(2245) ,
  \747GAT(219) ,
  \2657GAT(879) ,
  \3111GAT(1061) ,
  \894GAT(170) ,
  \4384GAT(1600) ,
  \2142GAT(624) ,
  \1413GAT(343) ,
  \1885GAT(509) ,
  \3244GAT(1115) ,
  \5410GAT(2040) ,
  \4583GAT(1671) ,
  \2656GAT(886) ,
  \918GAT(162) ,
  \3612GAT(1293) ,
  \978GAT(142) ,
  \1920GAT(554) ,
  \5422GAT(2035) ,
  \1327GAT(298) ,
  \3055GAT(1039) ,
  \2700GAT(904) ,
  \2046GAT(619) ,
  \4461GAT(1624) ,
  \2030GAT(578) ,
  \4048GAT(1455) ,
  \4554GAT(1680) ,
  \2823GAT(957) ,
  \4801GAT(1794) ,
  \3494GAT(1233) ,
  \3533GAT(1221) ,
  \5825GAT(2218) ,
  \2635GAT(848) ,
  \3331GAT(1162) ,
  \5705GAT(2176) ,
  \4642GAT(1716) ,
  \1053GAT(117) ,
  \5357GAT(2013) ,
  \5755GAT(2202) ,
  \1697GAT(458) ,
  \3830GAT(1385) ,
  \3049GAT(1041) ,
  \1600GAT(416) ,
  \1107GAT(99) ,
  \5831GAT(2215) ,
  \3923GAT(1410) ,
  \618GAT(262) ,
  \3361GAT(1151) ,
  \678GAT(242) ,
  \3221GAT(1124) ,
  \2712GAT(900) ,
  \5938GAT(2288) ,
  \2579GAT(828) ,
  \3902GAT(1419) ,
  \3505GAT(1244) ,
  \5214GAT(1971) ,
  \3628GAT(1289) ,
  \4172GAT(1495) ,
  \3658GAT(1278) ,
  \5573GAT(2120) ,
  \4956GAT(1870) ,
  \828GAT(192) ,
  \3127GAT(1054) ,
  \888GAT(172) ,
  \4851GAT(1806) ,
  \3739GAT(1329) ,
  \4090GAT(1478) ,
  \2655GAT(881) ,
  \4737GAT(1755) ,
  \4566GAT(1689) ,
  \2109GAT(634) ,
  \3860GAT(1377) ,
  \2346GAT(722) ,
  \5898GAT(2268) ,
  \4604GAT(1715) ,
  \2289GAT(711) ,
  \660GAT(248) ,
  \1726GAT(480) ,
  \2251GAT(690) ,
  \3310GAT(1137) ,
  \4793GAT(1783) ,
  \4290GAT(1564) ,
  \1884GAT(505) ,
  \3368GAT(1194) ,
  \6225GAT(2415) ,
  \3842GAT(1395) ,
  \3747GAT(1327) ,
  \1095GAT(103) ,
  \3322GAT(1130) ,
  \4524GAT(1688) ,
  \6211GAT(2407) ,
  \3931GAT(1418) ,
  \4357GAT(1612) ,
  \4173GAT(1537) ,
  \3699GAT(1296) ,
  \1987GAT(567) ,
  \5581GAT(2117) ,
  \3896GAT(1422) ,
  \1850GAT(530) ,
  \2654GAT(887) ,
  \4578GAT(1672) ,
  \3712GAT(1339) ,
  \4689GAT(1729) ,
  \5230GAT(1970) ,
  \5032GAT(1890) ,
  \2706GAT(902) ,
  \708GAT(232) ,
  \1698GAT(455) ,
  \1407GAT(345) ,
  \2650GAT(841) ,
  \4237GAT(1519) ,
  \3562GAT(1271) ,
  \2518GAT(800) ,
  \3157GAT(1101) ,
  \4058GAT(1489) ,
  \2999GAT(1014) ,
  \3193GAT(1075) ,
  \756GAT(216) ,
  \2227GAT(698) ,
  \1029GAT(125) ,
  \4456GAT(1625) ,
  \3280GAT(1144) ,
  \1664GAT(430) ,
  \1089GAT(105) ,
  \2539GAT(786) ,
  \3821GAT(1344) ,
  \3813GAT(1347) ,
  \2878GAT(982) ,
  \4220GAT(1535) ,
  \1699GAT(456) ,
  \4414GAT(1638) ,
  \2166GAT(674) ,
  \585GAT(273) ,
  \1410GAT(344) ,
  \3004GAT(1019) ,
  \4932GAT(1825) ,
  \2392GAT(751) ,
  \2164GAT(669) ,
  \4031GAT(1450) ,
  \2434GAT(777) ,
  \975GAT(143) ,
  \4802GAT(1781) ,
  \6286GAT(2446) ,
  \2149GAT(678) ,
  \5941GAT(2287) ,
  \3233GAT(1118) ,
  \1923GAT(553) ,
  \4833GAT(1817) ,
  \5409GAT(2051) ,
  \4964GAT(1868) ,
  \3404GAT(1180) ,
  \4078GAT(1492) ,
  \3334GAT(1171) ,
  \5866GAT(2254) ,
  \5184GAT(1975) ,
  \2368GAT(761) ,
  \6231GAT(2417) ,
  \5092GAT(1911) ,
  \3070GAT(1035) ,
  \6102GAT(2349) ,
  \4858GAT(1805) ,
  \6002GAT(2297) ,
  \3180GAT(1079) ,
  \6124GAT(2367) ,
  \5073GAT(1917) ,
  \6090GAT(2354) ,
  \4507GAT(1652) ,
  \2990GAT(1030) ,
  \2757GAT(922) ,
  \6040GAT(2335) ,
  \3062GAT(1038) ,
  \675GAT(243) ,
  \2831GAT(940) ,
  \5933GAT(2289) ,
  \5683GAT(2182) ,
  \1811GAT(488) ,
  \5226GAT(1957) ,
  \4899GAT(1836) ,
  \6207GAT(2404) ,
  \4854GAT(1815) ,
  \1323GAT(299) ,
  \4327GAT(1581) ,
  \3040GAT(1046) ,
  \3653GAT(1279) ,
  \3942GAT(1404) ,
  \6130GAT(2364) ,
  \3224GAT(1123) ,
  \900GAT(168) ,
  \1603GAT(415) ,
  \3141GAT(1108) ,
  \4232GAT(1520) ,
  \732GAT(224) ,
  \3254GAT(1111) ,
  \3260GAT(1109) ,
  \4953GAT(1871) ,
  \1779GAT(496) ,
  \5467GAT(2062) ,
  \1404GAT(346) ,
  \4007GAT(1461) ,
  \4106GAT(1472) ,
  \1889GAT(503) ,
  \4411GAT(1640) ,
  \6069GAT(2345) ,
  \2977GAT(986) ,
  \1648GAT(434) ,
  \2744GAT(889) ,
  \2837GAT(950) ,
  \1652GAT(433) ,
  \2422GAT(780) ,
  \4717GAT(1771) ,
  \3845GAT(1381) ,
  \2064GAT(613) ,
  \5972GAT(2308) ,
  \5327GAT(2034) ,
  \4423GAT(1645) ,
  \5455GAT(2079) ,
  \5005GAT(1902) ,
  \2508GAT(806) ,
  \2165GAT(676) ,
  \6261GAT(2432) ,
  \5553GAT(2132) ,
  \4779GAT(1789) ,
  \3392GAT(1192) ,
  \903GAT(167) ,
  \3389GAT(1184) ,
  \3797GAT(1352) ,
  \2761GAT(921) ,
  \2105GAT(635) ,
  \3664GAT(1313) ,
  \5389GAT(2047) ,
  \3735GAT(1340) ,
  \3003GAT(1011) ,
  \3007GAT(1009) ,
  \1839GAT(532) ,
  \5595GAT(2128) ,
  \3727GAT(1332) ,
  \3757GAT(1323) ,
  \2576GAT(830) ,
  \1486GAT(352) ,
  \1836GAT(537) ,
  \5043GAT(1887) ,
  \6236GAT(2421) ,
  \3099GAT(1064) ,
  \3670GAT(1308) ,
  \3323GAT(1170) ,
  \4775GAT(1798) ,
  \4563GAT(1676) ,
  \5056GAT(1882) ,
  \588GAT(272) ,
  \2285GAT(712) ,
  \1807GAT(489) ,
  \4028GAT(1451) ,
  \2627GAT(850) ,
  \2659GAT(877) ,
  \5780GAT(2193) ,
  \4339GAT(1576) ,
  \3602GAT(1255) ,
  \3198GAT(1074) ,
  \825GAT(193) ,
  \4541GAT(1694) ,
  \4217GAT(1524) ,
  \2169GAT(666) ,
  \2313GAT(705) ,
  \5968GAT(2277) ,
  \4194GAT(1543) ,
  \3702GAT(1305) ,
  \3911GAT(1415) ,
  \3353GAT(1153) ,
  \3115GAT(1060) ,
  \3852GAT(1391) ,
  \5787GAT(2230) ,
  \3236GAT(1117) ,
  \2658GAT(885) ,
  \4725GAT(1760) ,
  \4140GAT(1505) ,
  \3894GAT(1367) ,
  \855GAT(183) ,
  \981GAT(141) ,
  \4758GAT(1748) ,
  \2975GAT(987) ,
  \5064GAT(1880) ,
  \1098GAT(102) ,
  \4453GAT(1626) ,
  \4362GAT(1618) ,
  \2709GAT(901) ,
  \5365GAT(2011) ,
  \4229GAT(1521) ,
  \1729GAT(479) ,
  \2438GAT(776) ,
  \1059GAT(115) ,
  \4814GAT(1776) ,
  \5106GAT(1907) ,
  \882GAT(174) ,
  \5315GAT(2027) ,
  \4912GAT(1833) ,
  \4500GAT(1653) ,
  \705GAT(233) ,
  \5633GAT(2160) ,
  \3581GAT(1262) ,
  \3160GAT(1085) ,
  \2478GAT(822) ,
  \2532GAT(793) ,
  \2921GAT(966) ,
  \2170GAT(673) ,
  \2374GAT(759) ,
  \2549GAT(839) ,
  \3636GAT(1284) ,
  \6097GAT(2350) ,
  \4251GAT(1566) ,
  \3989GAT(1428) ,
  \5151GAT(1950) ,
  \6035GAT(2333) ,
  \5979GAT(2305) ,
  \4821GAT(1820) ,
  \4344GAT(1585) ,
  \2533GAT(791) ,
  \1859GAT(520) ,
  \6019GAT(2321) ,
  \6057GAT(2327) ,
  \2171GAT(671) ,
  \4089GAT(1477) ,
  \2922GAT(972) ,
  \2067GAT(612) ,
  \4920GAT(1830) ,
  \1834GAT(535) ,
  \3172GAT(1093) ,
  \5383GAT(2054) ,
  \3151GAT(1104) ,
  \993GAT(137) ,
  \4155GAT(1508) ,
  \1835GAT(539) ,
  \5380GAT(2049) ,
  \783GAT(207) ,
  \1775GAT(497) ,
  \2001GAT(562) ,
  \4784GAT(1787) ,
  \3980GAT(1435) ,
  \4643GAT(1702) ,
  \1644GAT(435) ,
  \5796GAT(2228) ,
  \4285GAT(1553) ,
  \4968GAT(1878) ,
  \4011GAT(1459) ,
  \3197GAT(1073) ,
  \2145GAT(623) ,
  \3831GAT(1400) ,
  \3685GAT(1302) ,
  \3326GAT(1175) ,
  \1026GAT(126) ,
  \693GAT(237) ,
  \669GAT(245) ,
  \3272GAT(1146) ,
  \5564GAT(2122) ,
  \990GAT(138) ,
  \4536GAT(1696) ,
  \4361GAT(1608) ,
  \5053GAT(1883) ,
  \4712GAT(1764) ,
  \4666GAT(1737) ,
  \5339GAT(2019) ,
  \6266GAT(2436) ,
  \2000GAT(564) ,
  \1419GAT(341) ,
  \3441GAT(1210) ,
  \6191GAT(2397) ,
  \3514GAT(1227) ,
  \2684GAT(861) ,
  \3074GAT(1033) ,
  \2923GAT(965) ,
  \912GAT(164) ,
  \690GAT(238) ,
  \5176GAT(1977) ,
  \3356GAT(1152) ,
  \3772GAT(1362) ,
  \1632GAT(438) ,
  \5697GAT(2178) ,
  \5628GAT(2150) ,
  \5352GAT(2015) ,
  \6167GAT(2384) ,
  \2052GAT(617) ,
  \4697GAT(1738) ,
  \1691GAT(464) ,
  \5913GAT(2263) ,
  \1609GAT(413) ,
  \2317GAT(702) ,
  \5296GAT(1981) ,
  \2377GAT(758) ,
  \2531GAT(788) ,
  \3540GAT(1220) ,
  \3465GAT(1199) ,
  \3340GAT(1165) ,
  \3748GAT(1325) ,
  \4319GAT(1588) ,
  \5180GAT(1976) ,
  \5277GAT(1987) ,
  \4474GAT(1665) ,
  \612GAT(264) ,
  \738GAT(222) ,
  \3930GAT(1409) ,
  \4813GAT(1778) ,
  \[0] ,
  \3825GAT(1387) ,
  \5654GAT(2158) ,
  \[1] ,
  \3873GAT(1374) ,
  \5980GAT(2306) ,
  \4551GAT(1690) ,
  \2687GAT(860) ,
  \[2] ,
  \5413GAT(2039) ,
  \[3] ,
  \3780GAT(1360) ,
  \6155GAT(2380) ,
  \[4] ,
  \3855GAT(1378) ,
  \822GAT(194) ,
  \[5] ,
  \2938GAT(999) ,
  \5679GAT(2184) ,
  \[6] ,
  \3230GAT(1120) ,
  \2976GAT(990) ,
  \3317GAT(1131) ,
  \[7] ,
  \3484GAT(1238) ,
  \5425GAT(2077) ,
  \[8] ,
  \4746GAT(1753) ,
  \4016GAT(1466) ,
  \[9] ,
  \4150GAT(1501) ,
  \2989GAT(1024) ,
  \720GAT(228) ,
  \2402GAT(749) ,
  \3016GAT(1007) ,
  \3662GAT(1315) ,
  \1690GAT(463) ,
  \780GAT(208) ,
  \1528GAT(393) ,
  \5155GAT(1936) ,
  \3300GAT(1136) ,
  \3947GAT(1443) ,
  \4870GAT(1800) ,
  \1855GAT(527) ,
  \5204GAT(1963) ,
  \1056GAT(116) ,
  \2476GAT(816) ,
  \5167GAT(1931) ,
  \5097GAT(1923) ,
  \666GAT(246) ,
  \5956GAT(2282) ,
  \5388GAT(2053) ,
  \3881GAT(1371) ,
  \1840GAT(536) ,
  \5239GAT(1999) ,
  \5671GAT(2137) ,
  \924GAT(160) ,
  \5066GAT(1929) ,
  \2653GAT(883) ,
  \858GAT(182) ,
  \2994GAT(1028) ,
  \2887GAT(979) ,
  \3899GAT(1421) ,
  \6020GAT(2317) ,
  \582GAT(274) ,
  \6187GAT(2394) ,
  \3837GAT(1397) ,
  \5459GAT(2065) ,
  \3977GAT(1431) ,
  \2506GAT(798) ,
  \6216GAT(2411) ,
  \5507GAT(2094) ,
  \5070GAT(1927) ,
  \5613GAT(2163) ,
  \2477GAT(823) ,
  \3715GAT(1338) ,
  \3985GAT(1434) ,
  \4077GAT(1482) ,
  \2838GAT(948) ,
  \5404GAT(2052) ,
  \723GAT(227) ,
  \1723GAT(481) ,
  \1693GAT(462) ,
  \4889GAT(1840) ,
  \1771GAT(498) ,
  \6106GAT(2361) ,
  \4364GAT(1617) ,
  \5516GAT(2092) ,
  \6175GAT(2390) ,
  \1494GAT(350) ,
  \6145GAT(2375) ,
  \5621GAT(2153) ,
  \2561GAT(835) ,
  \1367GAT(288) ,
  \5658GAT(2141) ,
  \1891GAT(504) ,
  \645GAT(253) ,
  \891GAT(171) ,
  \4943GAT(1822) ,
  \3998GAT(1424) ,
  \3043GAT(1044) ,
  \1416GAT(342) ,
  \4486GAT(1659) ,
  \1955GAT(575) ,
  \1692GAT(461) ,
  \5082GAT(1915) ,
  \1890GAT(506) ,
  \1372GAT(331) ,
  \927GAT(159) ,
  \5235GAT(1969) ,
  \3028GAT(1050) ,
  \6001GAT(2299) ,
  \6129GAT(2366) ,
  \1841GAT(534) ,
  \5946GAT(2286) ,
  \1854GAT(523) ,
  \2836GAT(937) ,
  \4179GAT(1549) ,
  \4265GAT(1561) ,
  \4098GAT(1475) ,
  \786GAT(206) ,
  \2019GAT(592) ,
  \2211GAT(647) ,
  \1032GAT(124) ,
  \4894GAT(1838) ,
  \5934GAT(2294) ,
  \735GAT(223) ,
  \4654GAT(1745) ,
  \3868GAT(1375) ,
  \3590GAT(1260) ,
  \4692GAT(1739) ,
  \1905GAT(559) ,
  \2362GAT(763) ,
  \6195GAT(2400) ,
  \2769GAT(919) ,
  \1983GAT(568) ,
  \4449GAT(1639) ,
  \2743GAT(888) ,
  \2896GAT(976) ,
  \3709GAT(1341) ,
  \2971GAT(991) ,
  \4310GAT(1590) ,
  \2133GAT(628) ,
  \3624GAT(1290) ,
  \3935GAT(1407) ,
  \1373GAT(330) ,
  \4198GAT(1530) ,
  \6277GAT(2439) ,
  \3409GAT(1179) ,
  \2993GAT(1020) ,
  \954GAT(150) ,
  \5168GAT(1932) ,
  \3119GAT(1057) ,
  \1556GAT(376) ,
  \2884GAT(980) ,
  \1938GAT(548) ,
  \1897GAT(501) ,
  \5026GAT(1897) ,
  \2210GAT(649) ,
  \3421GAT(1215) ,
  \4085GAT(1479) ,
  \5038GAT(1888) ,
  \1680GAT(426) ,
  \3176GAT(1092) ,
  \2930GAT(1001) ,
  \5959GAT(2281) ,
  \5975GAT(2307) ,
  \2430GAT(778) ,
  \654GAT(250) ,
  \5440GAT(2071) ,
  \5400GAT(2044) ,
  \3433GAT(1212) ,
  \1856GAT(525) ,
  \576GAT(276) ,
  \3339GAT(1157) ,
  \4570GAT(1675) ,
  \1557GAT(377) ,
  \3520GAT(1236) ,
  \2545GAT(783) ,
  \4386GAT(1599) ,
  \1606GAT(414) ,
  \5651GAT(2142) ,
  \5450GAT(2067) ,
  \4934GAT(1824) ,
  \3332GAT(1172) ,
  \3288GAT(1142) ,
  \4348GAT(1574) ,
  \1513GAT(402) ,
  \5322GAT(2024) ,
  \3677GAT(1314) ,
  \3545GAT(1218) ,
  \1687GAT(468) ,
  \3669GAT(1319) ,
  \5540GAT(2135) ,
  \2093GAT(638) ,
  \648GAT(252) ,
  \3245GAT(1113) ,
  \5706GAT(2174) ,
  \3736GAT(1330) ,
  \1720GAT(482) ,
  \2319GAT(701) ,
  \2160GAT(679) ,
  \5360GAT(2012) ,
  \4972GAT(1865) ,
  \4460GAT(1623) ,
  \4373GAT(1615) ,
  \3532GAT(1223) ,
  \4582GAT(1670) ,
  \3449GAT(1208) ,
  \3760GAT(1365) ,
  \6138GAT(2372) ,
  \3350GAT(1154) ,
  \4226GAT(1522) ,
  \4881GAT(1853) ,
  \4891GAT(1849) ,
  \2832GAT(953) ,
  \4616GAT(1724) ,
  \1062GAT(114) ,
  \2544GAT(785) ,
  \1302GAT(34) ,
  \5624GAT(2152) ,
  \837GAT(189) ,
  \3806GAT(1348) ,
  \2454GAT(772) ,
  \1861GAT(522) ,
  \1512GAT(404) ,
  \6201GAT(2402) ,
  \3922GAT(1412) ,
  \1995GAT(565) ,
  \4980GAT(1862) ,
  \4726GAT(1769) ,
  \1371GAT(332) ,
  \3861GAT(1388) ,
  \2014GAT(593) ,
  \1422GAT(340) ,
  \1686GAT(467) ,
  \3586GAT(1270) ,
  \1308GAT(32) ,
  \5421GAT(2037) ,
  \4260GAT(1562) ,
  \2833GAT(951) ,
  \3311GAT(1133) ,
  \3252GAT(1112) ,
  \3574GAT(1265) ,
  \1717GAT(483) ,
  \6058GAT(2325) ,
  \4184GAT(1547) ,
  \1908GAT(558) ,
  \2015GAT(596) ,
  \1713GAT(442) ,
  \2058GAT(615) ,
  \5616GAT(2154) ,
  \1305GAT(33) ,
  \5535GAT(2086) ,
  \1656GAT(432) ,
  \3751GAT(1335) ,
  \1959GAT(574) ,
  \2697GAT(905) ,
  \2037GAT(622) ,
  \2161GAT(677) ,
  \4356GAT(1621) ,
  \987GAT(139) ,
  \4521GAT(1646) ,
  \4022GAT(1464) ,
  \1860GAT(524) ,
  \5429GAT(2074) ,
  \4171GAT(1494) ,
  \4478GAT(1664) ,
  \4466GAT(1667) ,
  \4408GAT(1642) ,
  \2318GAT(704) ,
  \5023GAT(1892) ,
  \1935GAT(549) ,
  \2690GAT(859) ,
  \2765GAT(920) ,
  \5830GAT(2217) ,
  \4100GAT(1474) ,
  \1526GAT(394) ,
  \4850GAT(1808) ,
  \1511GAT(403) ,
  \1482GAT(353) ,
  \2998GAT(1025) ,
  \1712GAT(441) ,
  \1803GAT(490) ,
  \4539GAT(1684) ,
  \852GAT(184) ,
  \4242GAT(1570) ,
  \1849GAT(526) ,
  \4193GAT(1531) ,
  \3647GAT(1281) ,
  \5163GAT(1933) ,
  \2446GAT(774) ,
  \1689GAT(466) ,
  \3396GAT(1183) ,
  \3553GAT(1274) ,
  \5725GAT(2168) ,
  \4628GAT(1707) ,
  \4557GAT(1679) ,
  \5121GAT(1947) ,
  \1894GAT(502) ,
  \3678GAT(1303) ,
  \1932GAT(550) ,
  \2623GAT(851) ,
  \3187GAT(1084) ,
  \3698GAT(1298) ,
  \3470GAT(1206) ,
  \5569GAT(2131) ,
  \6036GAT(2336) ,
  \2843GAT(945) ,
  \4993GAT(1858) ,
  \2293GAT(710) ,
  \5215GAT(1960) ,
  \5200GAT(1965) ,
  \5130GAT(1952) ,
  \2016GAT(591) ,
  \3504GAT(1231) ,
  \1527GAT(395) ,
  \4238GAT(1517) ,
  \4499GAT(1655) ,
  \5748GAT(2210) ,
  \2842GAT(947) ,
  \6285GAT(2445) ,
  \3377GAT(1189) ,
  \5819GAT(2220) ,
  \4429GAT(1634) ,
  \4417GAT(1637) ,
  \3479GAT(1241) ,
  \5031GAT(1896) ,
  \5392GAT(2046) ,
  \3721GAT(1336) ,
  \4535GAT(1697) ,
  \5877GAT(2239) ,
  \2018GAT(589) ,
  \5528GAT(2087) ,
  \1711GAT(444) ,
  \3595GAT(1258) ,
  \5892GAT(2270) ,
  \5276GAT(2000) ,
  \999GAT(135) ,
  \5102GAT(1922) ,
  \4146GAT(1503) ,
  \4380GAT(1602) ,
  \4269GAT(1571) ,
  \1517GAT(401) ,
  \729GAT(225) ,
  \789GAT(205) ,
  \4257GAT(1563) ,
  \4368GAT(1616) ,
  \5093GAT(1912) ,
  \3800GAT(1351) ,
  \5113GAT(1904) ,
  \1688GAT(465) ,
  \996GAT(136) ,
  \5227GAT(1955) ,
  \2739GAT(890) ,
  \6103GAT(2347) ,
  \2017GAT(594) ,
  \5694GAT(2179) ,
  \2694GAT(906) ,
  \6091GAT(2352) ,
  \2156GAT(680) ,
  \5301GAT(1979) ,
  \5852GAT(2248) ,
  \3031GAT(1049) ,
  \699GAT(235) ,
  \4687GAT(1730) ,
  \4094GAT(1487) ,
  \1521GAT(397) ,
  \3616GAT(1292) ,
  \984GAT(140) ,
  \5718GAT(2171) ,
  \4006GAT(1471) ,
  \1038GAT(122) ,
  \2010GAT(597) ,
  \1710GAT(443) ,
  \2458GAT(771) ,
  \2371GAT(760) ,
  \1537GAT(389) ,
  \5209GAT(1972) ,
  \696GAT(236) ,
  \5659GAT(2157) ,
  \1516GAT(400) ,
  \1454GAT(360) ,
  \3882GAT(1380) ,
  \2615GAT(853) ,
  \4658GAT(1744) ,
  \5333GAT(2021) ,
  \3002GAT(1021) ,
  \3142GAT(1107) ,
  \3314GAT(1132) ,
  \5118GAT(1948) ,
  \4872GAT(1799) ,
  \1947GAT(577) ,
  \6156GAT(2381) ,
  \3474GAT(1197) ,
  \2926GAT(1002) ,
  \2155GAT(681) ,
  \4328GAT(1586) ,
  \606GAT(266) ,
  \5134GAT(1943) ,
  \6257GAT(2429) ,
  \4027GAT(1462) ,
  \1522GAT(398) ,
  \1999GAT(563) ,
  \5473GAT(2059) ,
  \6206GAT(2406) ,
  \3665GAT(1321) ,
  \2154GAT(675) ,
  \867GAT(179) ,
  \2139GAT(625) ,
  \834GAT(190) ,
  \6247GAT(2424) ,
  \3475GAT(1205) ,
  \1558GAT(375) ,
  \5585GAT(2115) ,
  \5515GAT(2106) ,
  \3027GAT(1004) ,
  \3693GAT(1299) ,
  \3058GAT(1045) ,
  \3133GAT(1051) ,
  \4019GAT(1453) ,
  \2841GAT(935) ,
  \5810GAT(2222) ,
  \5801GAT(2226) ,
  \1536GAT(388) ,
  \2138GAT(627) ,
  \3794GAT(1353) ,
  \2853GAT(939) ,
  \5743GAT(2211) ,
  \3846GAT(1394) ,
  \2055GAT(616) ,
  \1379GAT(324) ,
  \2934GAT(1000) ,
  \1941GAT(547) ,
  \3690GAT(1300) ,
  \4052GAT(1491) ,
  \2899GAT(975) ,
  \4353GAT(1614) ,
  \4733GAT(1757) ,
  \5596GAT(2112) ,
  \3724GAT(1334) ,
  \3268GAT(1147) ,
  \3413GAT(1185) ,
  \4714GAT(1763) ,
  \5042GAT(1886) ,
  \6235GAT(2420) ,
  \2852GAT(941) ,
  \1523GAT(396) ,
  \5379GAT(2055) ,
  \4839GAT(1811) ,
  \3335GAT(1159) ,
  \5865GAT(2244) ,
  \4444GAT(1641) ,
  \5495GAT(2099) ,
  \771GAT(211) ,
  \5527GAT(2089) ,
  \3284GAT(1143) ,
  \1846GAT(531) ,
  \4884GAT(1841) ,
  \4562GAT(1678) ,
  \6176GAT(2391) ,
  \5945GAT(2285) ,
  \2997GAT(1016) ,
  \5489GAT(2109) ,
  \4540GAT(1695) ,
  \5114GAT(1905) ,
  \1636GAT(437) ,
  \609GAT(265) ,
  \5781GAT(2194) ,
  \3481GAT(1253) ,
  \3491GAT(1249) ,
  \1068GAT(112) ,
  \4195GAT(1542) ,
  \4701GAT(1726) ,
  \5700GAT(2177) ,
  \1378GAT(325) ,
  \2012GAT(595) ,
  \1844GAT(529) ,
  \2297GAT(709) ,
  \5094GAT(1910) ,
  \2407GAT(747) ,
  \3445GAT(1209) ,
  \2683GAT(866) ,
  \6161GAT(2382) ,
  \1458GAT(359) ,
  \4503GAT(1661) ,
  \921GAT(161) ,
  \4759GAT(1749) ,
  \4890GAT(1850) ,
  \1035GAT(123) ,
  \579GAT(275) ,
  \2013GAT(598) ,
  \2567GAT(833) ,
  \6146GAT(2376) ,
  \5786GAT(2237) ,
  \5364GAT(2010) ,
  \6134GAT(2371) ,
  \2205GAT(652) ,
  \5857GAT(2247) ,
  \1498GAT(349) ,
  \5988GAT(2303) ,
  \5146GAT(1938) ,
  \5663GAT(2139) ,
  \4911GAT(1832) ,
  \6009GAT(2320) ,
  \2322GAT(703) ,
  \864GAT(180) ,
  \6094GAT(2351) ,
  \5773GAT(2196) ,
  \4584GAT(1669) ,
  \3208GAT(1070) ,
  \3657GAT(1277) ,
  \6044GAT(2331) ,
  \4808GAT(1779) ,
  \2206GAT(650) ,
  \4188GAT(1532) ,
  \4667GAT(1742) ,
  \2564GAT(834) ,
  \3938GAT(1406) ,
  \4763GAT(1793) ,
  \4010GAT(1469) ,
  \3742GAT(1328) ,
  \2773GAT(918) ,
  \5962GAT(2280) ,
  \5256GAT(2002) ,
  \4323GAT(1587) ,
  \3641GAT(1286) ,
  \4274GAT(1569) ,
  \3152GAT(1103) ,
  \3175GAT(1081) ,
  \2851GAT(933) ,
  \3365GAT(1195) ,
  \6181GAT(2392) ,
  \5834GAT(2253) ,
  \4713GAT(1773) ,
  \6118GAT(2357) ,
  \4632GAT(1705) ,
  \2682GAT(862) ,
  \4986GAT(1859) ,
  \2619GAT(852) ,
  \2736GAT(891) ,
  \3963GAT(1439) ,
  \3171GAT(1095) ,
  \2217GAT(643) ,
  \1951GAT(576) ,
  \5387GAT(2048) ,
  \5443GAT(2070) ,
  \5292GAT(1998) ,
  \5950GAT(2292) ,
  \1490GAT(351) ,
  \4738GAT(1756) ,
  \1591GAT(419) ,
  \3348GAT(1155) ,
  \4937GAT(1839) ,
  \1363GAT(289) ,
  \5431GAT(2073) ,
  \1375GAT(328) ,
  \3971GAT(1437) ,
  \6265GAT(2435) ,
  \3383GAT(1187) ,
  \3548GAT(1217) ,
  \5602GAT(2110) ,
  \3292GAT(1141) ,
  \4286GAT(1554) ,
  \2552GAT(838) ,
  \2194GAT(651) ,
  \4372GAT(1605) ,
  \2121GAT(631) ,
  \1428GAT(338) ,
  \2607GAT(855) ,
  \5565GAT(2123) ,
  \4959GAT(1869) ,
  \4721GAT(1770) ,
  \3674GAT(1306) ,
  \1869GAT(514) ,
  \2675GAT(863) ,
  \5578GAT(2118) ,
  \4204GAT(1539) ,
  \2543GAT(784) ,
  \2881GAT(981) ,
  \4047GAT(1445) ,
  \1845GAT(533) ,
  \4675GAT(1735) ,
  \4401GAT(1595) ,
  \5370GAT(2057) ,
  \5768GAT(2198) ,
  \5493GAT(2100) ,
  \5088GAT(1913) ,
  \5912GAT(2272) ,
  \2404GAT(748) ,
  \567GAT(279) ,
  \726GAT(226) ,
  \3788GAT(1358) ,
  \4039GAT(1448) ,
  \2195GAT(658) ,
  \5246GAT(2006) ,
  \3531GAT(1222) ,
  \1374GAT(329) ,
  \957GAT(149) ,
  \642GAT(254) ,
  \4138GAT(1506) ,
  \831GAT(191) ,
  \5557GAT(2125) ,
  \5714GAT(2188) ,
  \6111GAT(2360) ,
  \4134GAT(1510) ,
  \3686GAT(1310) ,
  \3862GAT(1386) ,
  \3992GAT(1427) ,
  \2159GAT(672) ,
  \4190GAT(1544) ,
  \3856GAT(1390) ,
  \5629GAT(2151) ,
  \3455GAT(1203) ,
  \2386GAT(755) ,
  \4751GAT(1751) ,
  \3889GAT(1368) ,
  \3638GAT(1283) ,
  \5981GAT(2304) ,
  \5776GAT(2195) ,
  \2137GAT(626) ,
  \1685GAT(425) ,
  \1041GAT(121) ,
  \2403GAT(752) ,
  \3663GAT(1322) ,
  \3362GAT(1149) ,
  \5903GAT(2267) ,
  \5769GAT(2208) ,
  \4747GAT(1765) ,
  \657GAT(249) ,
  \1767GAT(499) ,
  \5156GAT(1949) ,
  \2806GAT(955) ,
  \6271GAT(2437) ,
  \2988GAT(1031) ,
  \3840GAT(1383) ,
  \2807GAT(964) ,
  \4103GAT(1473) ,
  \3327GAT(1166) ,
  \2196GAT(656) ,
  \5666GAT(2138) ,
  \1377GAT(326) ,
  \4550GAT(1691) ,
  \2893GAT(977) ,
  \5172GAT(1945) ,
  \2674GAT(870) ,
  \5789GAT(2229) ,
  \3730GAT(1342) ,
  \3207GAT(1078) ,
  \4534GAT(1685) ,
  \4151GAT(1502) ,
  \4611GAT(1712) ,
  \2332GAT(736) ,
  \1553GAT(378) ,
  \5630GAT(2149) ,
  \951GAT(151) ,
  \4662GAT(1743) ,
  \1538GAT(387) ,
  \1967GAT(572) ,
  \1065GAT(113) ,
  \6227GAT(2414) ,
  \4355GAT(1613) ,
  \5067GAT(1920) ,
  \4164GAT(1497) ,
  \5590GAT(2129) ,
  \2214GAT(644) ,
  \1747GAT(473) ,
  \4183GAT(1534) ,
  \3121GAT(1056) ,
  \1684GAT(424) ,
  \3792GAT(1354) ,
  \5160GAT(1934) ,
  \2333GAT(741) ,
  \4625GAT(1708) ,
  \1864GAT(517) ,
  \3429GAT(1213) ,
  \3301GAT(1139) ,
  \5798GAT(2227) ,
  \1251GAT(51) ,
  \1431GAT(337) ,
  \1552GAT(380) ,
  \2731GAT(893) ,
  \5205GAT(1964) ,
  \1376GAT(327) ,
  \2097GAT(637) ,
  \2890GAT(978) ,
  \1254GAT(50) ,
  \4001GAT(1433) ,
  \4441GAT(1629) ,
  \3827GAT(1401) ,
  \1865GAT(521) ,
  \2803GAT(907) ,
  \651GAT(251) ,
  \2732GAT(897) ,
  \1991GAT(566) ,
  \5135GAT(1951) ,
  \3182GAT(1087) ,
  \2248GAT(691) ,
  \564GAT(280) ,
  \3276GAT(1145) ,
  \5739GAT(2212) ,
  \6215GAT(2410) ,
  \3328GAT(1174) ,
  \5244GAT(1997) ,
  \573GAT(277) ,
  \5142GAT(1940) ,
  \5891GAT(2274) ,
  \3598GAT(1257) ,
  \6107GAT(2363) ,
  \5408GAT(2041) ,
  \2450GAT(773) ,
  \3006GAT(1017) ,
  \3341GAT(1156) ,
  \1744GAT(474) ,
  \2329GAT(744) ,
  \3264GAT(1148) ,
  \5761GAT(2199) ,
  \936GAT(156) ,
  \4015GAT(1456) ,
  \5271GAT(2001) ,
  \3976GAT(1436) ,
  \1902GAT(560) ,
  \777GAT(209) ,
  \5955GAT(2291) ,
  \3386GAT(1186) ,
  \4281GAT(1555) ,
  \3951GAT(1442) ,
  \3243GAT(1114) ,
  \2027GAT(584) ,
  \4637GAT(1718) ,
  \4718GAT(1761) ,
  \4494GAT(1656) ,
  \3984GAT(1430) ,
  \4974GAT(1864) ,
  \4942GAT(1837) ,
  \5548GAT(2133) ,
  \3814GAT(1355) ,
  \5506GAT(2096) ,
  \4592GAT(1721) ,
  \5929GAT(2296) ,
  \5059GAT(1881) ,
  \3893GAT(1366) ,
  \6276GAT(2441) ,
  \4254GAT(1565) ,
  \3671GAT(1318) ,
  \2802GAT(909) ,
  \5760GAT(2201) ,
  \3490GAT(1250) ,
  \3083GAT(1068) ,
  \5822GAT(2219) ,
  \5967GAT(2279) ,
  \3768GAT(1363) ,
  \5752GAT(2203) ,
  \1914GAT(556) ,
  \2330GAT(738) ,
  \2328GAT(740) ,
  \570GAT(278) ,
  \5309GAT(2029) ,
  \636GAT(256) ,
  \4340GAT(1577) ,
  \1551GAT(379) ,
  \4199GAT(1541) ,
  \4515GAT(1649) ,
  \5001GAT(1855) ,
  \2026GAT(581) ,
  \2848GAT(942) ,
  \5574GAT(2130) ,
  \6000GAT(2298) ,
  \3877GAT(1382) ,
  \5649GAT(2143) ,
  \3218GAT(1125) ,
  \5236GAT(1953) ,
  \801GAT(201) ,
  \5904GAT(2265) ,
  \2389GAT(753) ,
  \2817GAT(960) ,
  \5071GAT(1918) ,
  \2082GAT(606) ,
  \3511GAT(1240) ,
  \1866GAT(519) ,
  \2678GAT(868) ,
  \5298GAT(1980) ,
  \3997GAT(1426) ,
  \6005GAT(2324) ,
  \1531GAT(391) ,
  \1381GAT(322) ,
  \2129GAT(629) ,
  \4904GAT(1835) ,
  \2442GAT(775) ,
  \2808GAT(963) ,
  \3706GAT(1343) ,
  \6080GAT(2338) ,
  \5318GAT(2026) ,
  \2733GAT(892) ,
  \4512GAT(1650) ,
  \963GAT(147) ,
  \711GAT(231) ,
  \2331GAT(743) ,
  \5103GAT(1908) ,
  \2801GAT(908) ,
  \2025GAT(586) ,
  \3776GAT(1361) ,
  \3344GAT(1163) ,
  \5017GAT(1899) ,
  \1425GAT(339) ,
  \3155GAT(1088) ,
  \2846GAT(934) ,
  \2847GAT(944) ,
  \6052GAT(2328) ,
  \2081GAT(609) ,
  \1359GAT(290) ,
  \2327GAT(745) ,
  \3022GAT(1005) ,
  \4009GAT(1460) ,
  \4995GAT(1857) ,
  \5461GAT(2064) ,
  \2464GAT(768) ,
  \2858GAT(936) ,
  \600GAT(268) ,
  \5139GAT(1941) ,
  \1799GAT(491) ,
  \1380GAT(323) ,
  \4349GAT(1584) ,
  \3371GAT(1193) ,
  \5692GAT(2180) ,
  \5846GAT(2250) ,
  \4742GAT(1767) ,
  \5169GAT(1930) ,
  \4482GAT(1663) ,
  \2992GAT(1029) ,
  \1566GAT(370) ,
  \5536GAT(2102) ,
  \5673GAT(2186) ,
  \2641GAT(843) ,
  \2818GAT(959) ,
  \5068GAT(1928) ,
  \6114GAT(2359) ,
  \1071GAT(111) ,
  \4470GAT(1666) ,
  \4448GAT(1628) ,
  \2958GAT(994) ,
  \4114GAT(1515) ,
  \3167GAT(1096) ,
  \2987GAT(1026) ,
  \1532GAT(392) ,
  \2640GAT(847) ,
  \4266GAT(1559) ,
  \4374GAT(1604) ,
  \3672GAT(1307) ,
  \3818GAT(1345) ,
  \5730GAT(2214) ,
  \1383GAT(320) ,
  \5638GAT(2159) ,
  \3666GAT(1311) ,
  \5660GAT(2140) ,
  \4561GAT(1677) ,
  \2080GAT(607) ,
  \5925GAT(2258) ,
  \4796GAT(1796) ;
assign
  \4248GAT(1567)  = ~\4189GAT(1545)  & ~\4188GAT(1532) ,
  \2326GAT(742)  = ~\2269GAT(716)  & ~\2224GAT(699) ,
  \2591GAT(829)  = ~\1230GAT(58)  & ~\2545GAT(783) ,
  \4126GAT(1512)  = ~\762GAT(214)  & ~\4064GAT(1486) ,
  \1870GAT(518)  = ~\981GAT(141)  & ~\1799GAT(491) ,
  \2467GAT(767)  = ~\2403GAT(752)  & ~\2402GAT(749) ,
  \603GAT(267)  = \341GAT(20)  & \18GAT(1) ,
  \1714GAT(440)  = ~\1685GAT(425)  & ~\1684GAT(424) ,
  \4278GAT(1556)  = ~\4225GAT(1533)  & ~\4224GAT(1523) ,
  \6177GAT(2389)  = ~\6171GAT(2387)  & ~\6076GAT(2340) ,
  \2024GAT(583)  = ~\1987GAT(567)  & ~\1932GAT(550) ,
  \4805GAT(1780)  = ~\4747GAT(1765)  & ~\4746GAT(1753) ,
  \1567GAT(371)  = ~\1122GAT(94)  & ~\1494GAT(350) ,
  \4215GAT(1525)  = ~\4146GAT(1503)  & ~\4082GAT(1480) ,
  \1533GAT(390)  = ~\1466GAT(357)  & ~\1331GAT(297) ,
  \4925GAT(1828)  = ~\4859GAT(1814)  & ~\4858GAT(1805) ,
  \6030GAT(2313)  = ~\5996GAT(2300)  & ~\5959GAT(2281) ,
  \2209GAT(645)  = ~\2133GAT(628)  & ~\2073GAT(608) ,
  \5617GAT(2162)  = ~\678GAT(242)  & ~\5548GAT(2133) ,
  \3145GAT(1094)  = ~\3083GAT(1068)  & ~\3031GAT(1049) ,
  \939GAT(155)  = \341GAT(20)  & \137GAT(8) ,
  \5785GAT(2231)  = ~\5730GAT(2214)  & ~\5673GAT(2186) ,
  \5374GAT(2056)  = ~\5251GAT(2004)  & ~\5315GAT(2027) ,
  \3784GAT(1359)  = ~\855GAT(183)  & ~\3724GAT(1334) ,
  \5254GAT(1994)  = ~\5188GAT(1974)  & ~\5127GAT(1944) ,
  \1621GAT(409)  = ~\1577GAT(365)  & ~\1576GAT(364) ,
  \4491GAT(1657)  = ~\4428GAT(1644)  & ~\4427GAT(1635) ,
  \1311GAT(302)  = ~\591GAT(271) ,
  \5428GAT(2083)  = ~\5246GAT(2006)  & ~\5370GAT(2057) ,
  \1450GAT(361)  = ~\594GAT(270)  & ~\1404GAT(346) ,
  \4963GAT(1867)  = ~\4907GAT(1834)  & ~\4842GAT(1810) ,
  \1382GAT(321)  = ~\1331GAT(297) ,
  \3496GAT(1247)  = ~\3429GAT(1213)  & ~\3276GAT(1145) ,
  \4901GAT(1845)  = ~\4833GAT(1817)  & ~\4662GAT(1743) ,
  \2611GAT(854)  = ~\2498GAT(812)  & ~\2561GAT(835) ,
  \4360GAT(1619)  = ~\4190GAT(1544)  & ~\4306GAT(1591) ,
  \4880GAT(1854)  = ~\576GAT(276)  & ~\4817GAT(1821) ,
  \6200GAT(2403)  = \[21] ,
  \2595GAT(858)  = ~\2478GAT(822)  & ~\2549GAT(839) ,
  \5052GAT(1894)  = ~\1158GAT(82)  & ~\4989GAT(1874) ,
  \1946GAT(546)  = ~\1821GAT(484)  & ~\1897GAT(501) ,
  \1917GAT(555)  = ~\1855GAT(527)  & ~\1854GAT(523) ,
  \1871GAT(516)  = ~\1799GAT(491)  & ~\1664GAT(430) ,
  \1672GAT(428)  = ~\1563GAT(372)  & ~\1615GAT(411) ,
  \639GAT(255)  = \273GAT(16)  & \35GAT(2) ,
  \3486GAT(1251)  = ~\3421GAT(1215)  & ~\3268GAT(1147) ,
  \762GAT(214)  = \426GAT(25)  & \69GAT(4) ,
  \3410GAT(1177)  = ~\3361GAT(1151)  & ~\3360GAT(1150) ,
  \3921GAT(1411)  = ~\3868GAT(1375)  & ~\3797GAT(1352) ,
  \960GAT(148)  = \460GAT(27)  & \137GAT(8) ,
  \2856GAT(931)  = ~\2785GAT(915)  & ~\2724GAT(894) ,
  \5266GAT(1990)  = ~\5200GAT(1965)  & ~\5139GAT(1941) ,
  \4320GAT(1582)  = ~\4265GAT(1561)  & ~\4264GAT(1560) ,
  \4208GAT(1528)  = ~\4139GAT(1509)  & ~\4138GAT(1506) ,
  \5606GAT(2156)  = ~\5540GAT(2135)  & ~\5480GAT(2105) ,
  \4350GAT(1573)  = ~\4290GAT(1564)  & ~\4106GAT(1472) ,
  \5420GAT(2036)  = ~\5360GAT(2012)  & ~\5301GAT(1979) ,
  \5770GAT(2197)  = ~\5709GAT(2189)  & ~\5522GAT(2090) ,
  \3333GAT(1160)  = ~\3284GAT(1143)  & ~\3227GAT(1122) ,
  \3577GAT(1264)  = ~\3521GAT(1234)  & ~\3524GAT(1225) ,
  \5684GAT(2183)  = ~\5554GAT(2126)  & ~\5624GAT(2152) ,
  \681GAT(241)  = \511GAT(30)  & \35GAT(2) ,
  \4185GAT(1546)  = ~\4118GAT(1514)  & ~\3955GAT(1441) ,
  \774GAT(210)  = \494GAT(29)  & \69GAT(4) ,
  \3850GAT(1379)  = ~\3780GAT(1360)  & ~\3721GAT(1336) ,
  \6251GAT(2427)  = ~\6247GAT(2424)  & ~\5879GAT(2238) ,
  \1347GAT(293)  = ~\1023GAT(127) ,
  \2151GAT(682)  = ~\2085GAT(640)  & ~\1947GAT(577) ,
  \3461GAT(1201)  = ~\3398GAT(1182)  & ~\3401GAT(1181) ,
  \3565GAT(1269)  = ~\3505GAT(1244)  & ~\3504GAT(1231) ,
  \5642GAT(2146)  = ~\5574GAT(2130)  & ~\5573GAT(2120) ,
  \3211GAT(1128)  = \[6] ,
  \5818GAT(2232)  = ~\1020GAT(128)  & ~\5764GAT(2209) ,
  \1002GAT(134)  = \426GAT(25)  & \154GAT(9) ,
  \2269GAT(716)  = ~\2151GAT(682)  & ~\2224GAT(699) ,
  \6241GAT(2422)  = ~\6237GAT(2419)  & ~\5925GAT(2258) ,
  \2946GAT(997)  = ~\2833GAT(951)  & ~\2893GAT(977) ,
  \6037GAT(2332)  = ~\6010GAT(2323)  & ~\6009GAT(2320) ,
  \3170GAT(1082)  = ~\3103GAT(1063)  & ~\3046GAT(1042) ,
  \2857GAT(938)  = ~\1038GAT(122)  & ~\2785GAT(915) ,
  \4520GAT(1648)  = ~\4395GAT(1597)  & ~\4456GAT(1625) ,
  \3646GAT(1285)  = ~\1095GAT(103)  & ~\3586GAT(1270) ,
  \5044GAT(1885)  = ~\4985GAT(1861)  & ~\4984GAT(1860) ,
  \2983GAT(984)  = ~\2923GAT(965)  & ~\1281GAT(41) ,
  \2245GAT(692)  = ~\2190GAT(661)  & ~\2189GAT(654) ,
  \846GAT(186)  = \358GAT(21)  & \103GAT(6) ,
  \5809GAT(2224)  = ~\5694GAT(2179)  & ~\5755GAT(2202) ,
  \5416GAT(2038)  = ~\5354GAT(2014)  & ~\5357GAT(2013) ,
  \1705GAT(450)  = ~\1553GAT(378)  & ~\1664GAT(430) ,
  \5251GAT(2004)  = ~\5184GAT(1975)  & ~\5013GAT(1900) ,
  \4727GAT(1759)  = ~\4671GAT(1741)  & ~\4494GAT(1656) ,
  \4428GAT(1644)  = ~\909GAT(165)  & ~\4368GAT(1616) ,
  \5747GAT(2205)  = ~\5688GAT(2191)  & ~\5630GAT(2149) ,
  \5676GAT(2185)  = ~\5617GAT(2162)  & ~\5616GAT(2154) ,
  \3253GAT(1119)  = ~\1188GAT(72)  & ~\3202GAT(1080) ,
  \3015GAT(1013)  = ~\1137GAT(89)  & ~\2971GAT(991) ,
  \4698GAT(1727)  = ~\4637GAT(1718)  & ~\4456GAT(1625) ,
  \3052GAT(1040)  = ~\3004GAT(1019)  & ~\3003GAT(1011) ,
  \2028GAT(579)  = ~\1995GAT(565)  & ~\1938GAT(548) ,
  \3552GAT(1275)  = \[7] ,
  \5726GAT(2169)  = ~\5596GAT(2112)  & ~\5666GAT(2138) ,
  \2200GAT(655)  = ~\1032GAT(124)  & ~\2125GAT(630) ,
  \5688GAT(2191)  = ~\825GAT(193)  & ~\5630GAT(2149) ,
  \4791GAT(1784)  = ~\4733GAT(1757)  & ~\4680GAT(1733) ,
  \5192GAT(1968)  = ~\5130GAT(1952)  & ~\5073GAT(1917) ,
  \2150GAT(683)  = ~\552GAT(284)  & ~\2085GAT(640) ,
  \5297GAT(1996)  = ~\1209GAT(65)  & ~\5230GAT(1970) ,
  \3832GAT(1399)  = ~\3764GAT(1364)  & ~\3608GAT(1294) ,
  \4650GAT(1746)  = ~\4531GAT(1698)  & ~\4595GAT(1720) ,
  \3019GAT(1006)  = ~\2976GAT(990)  & ~\2975GAT(987) ,
  \1945GAT(545)  = ~\1897GAT(501)  & ~\1269GAT(45) ,
  \5013GAT(1900)  = ~\4891GAT(1849)  & ~\4953GAT(1871) ,
  \1355GAT(291)  = ~\1119GAT(95) ,
  \4676GAT(1740)  = ~\960GAT(148)  & ~\4616GAT(1724) ,
  \2184GAT(657)  = ~\2113GAT(633)  & ~\2058GAT(615) ,
  \5030GAT(1891)  = ~\4968GAT(1878)  & ~\4913GAT(1831) ,
  \5022GAT(1898)  = ~\4901GAT(1845)  & ~\4959GAT(1869) ,
  \4359GAT(1610)  = ~\4306GAT(1591)  & ~\4251GAT(1566) ,
  \3425GAT(1214)  = ~\660GAT(248)  & ~\3371GAT(1193) ,
  \2011GAT(600)  = ~\1841GAT(534)  & ~\1959GAT(574) ,
  \5345GAT(2016)  = ~\5288GAT(1984)  & ~\5287GAT(1983) ,
  \861GAT(181)  = \443GAT(26)  & \103GAT(6) ,
  \4772GAT(1790)  = ~\4717GAT(1771)  & ~\4716GAT(1762) ,
  \804GAT(200)  = \392GAT(23)  & \86GAT(5) ,
  \4013GAT(1458)  = ~\3963GAT(1439)  & ~\3908GAT(1416) ,
  \3374GAT(1191)  = ~\3330GAT(1173)  & ~\3329GAT(1164) ,
  \4498GAT(1654)  = ~\4435GAT(1632)  & ~\4377GAT(1603) ,
  \6150GAT(2378)  = \[16] ,
  \3380GAT(1188)  = ~\3334GAT(1171)  & ~\3333GAT(1160) ,
  \5882GAT(2276)  = ~\585GAT(273)  & ~\5834GAT(2253) ,
  \6049GAT(2329)  = ~\6019GAT(2321)  & ~\6018GAT(2318) ,
  \4546GAT(1692)  = ~\4478GAT(1664)  & ~\4310GAT(1590) ,
  \3161GAT(1100)  = ~\753GAT(217)  & ~\3095GAT(1065) ,
  \3186GAT(1086)  = ~\993GAT(137)  & ~\3115GAT(1060) ,
  \2199GAT(648)  = ~\2125GAT(630)  & ~\2067GAT(612) ,
  \2029GAT(582)  = ~\1886GAT(507)  & ~\1995GAT(565) ,
  \1507GAT(407)  = ~\546GAT(286)  & ~\1446GAT(362) ,
  \4800GAT(1782)  = ~\4742GAT(1767)  & ~\4689GAT(1729) ,
  \3687GAT(1301)  = ~\3641GAT(1286)  & ~\3461GAT(1201) ,
  \4845GAT(1809)  = ~\4781GAT(1788)  & ~\4784GAT(1787) ,
  \3103GAT(1063)  = ~\849GAT(185)  & ~\3046GAT(1042) ,
  \2185GAT(664)  = ~\888GAT(172)  & ~\2113GAT(633) ,
  \2954GAT(995)  = ~\2843GAT(945)  & ~\2899GAT(975) ,
  \2201GAT(653)  = ~\2125GAT(630)  & ~\1987GAT(567) ,
  \1795GAT(492)  = ~\933GAT(157)  & ~\1741GAT(475) ,
  \3202GAT(1080)  = ~\1188GAT(72)  & ~\3133GAT(1051) ,
  \3437GAT(1211)  = ~\804GAT(200)  & ~\3380GAT(1188) ,
  \5332GAT(2033)  = ~\918GAT(162)  & ~\5271GAT(2001) ,
  \4064GAT(1486)  = ~\4014GAT(1467)  & ~\4013GAT(1458) ,
  \3536GAT(1230)  = ~\1143GAT(87)  & ~\3467GAT(1198) ,
  \5618GAT(2161)  = ~\5548GAT(2133)  & ~\5374GAT(2056) ,
  \2558GAT(836)  = ~\2497GAT(814)  & ~\2496GAT(804) ,
  \1568GAT(369)  = ~\1494GAT(350)  & ~\1359GAT(290) ,
  \4922GAT(1829)  = ~\4854GAT(1815)  & ~\4683GAT(1732) ,
  \6256GAT(2431)  = ~\6247GAT(2424)  & ~\6251GAT(2427) ,
  \5472GAT(2061)  = ~\5354GAT(2014)  & ~\5416GAT(2038) ,
  \3524GAT(1225)  = ~\3454GAT(1207)  & ~\3453GAT(1204) ,
  \2089GAT(639)  = ~\600GAT(268)  & ~\2040GAT(621) ,
  \3087GAT(1067)  = ~\657GAT(249)  & ~\3034GAT(1048) ,
  \4332GAT(1579)  = ~\4274GAT(1569)  & ~\4273GAT(1558) ,
  \3324GAT(1176)  = ~\3142GAT(1107)  & ~\3264GAT(1148) ,
  \4082GAT(1480)  = ~\4027GAT(1462)  & ~\4026GAT(1452) ,
  \4273GAT(1558)  = ~\4220GAT(1535)  & ~\4152GAT(1500) ,
  \4780GAT(1797)  = ~\864GAT(180)  & ~\4721GAT(1770) ,
  \5241GAT(2008)  = ~\5176GAT(1977)  & ~\5005GAT(1902) ,
  \2266GAT(684)  = ~\2222GAT(642)  & ~\2221GAT(641) ,
  \5544GAT(2134)  = ~\630GAT(258)  & ~\5483GAT(2103) ,
  \3926GAT(1420)  = ~\1050GAT(118)  & ~\3874GAT(1372) ,
  \3046GAT(1042)  = ~\3000GAT(1023)  & ~\2999GAT(1014) ,
  \4646GAT(1747)  = ~\4526GAT(1700)  & ~\4592GAT(1721) ,
  \2516GAT(792)  = ~\2446GAT(774)  & ~\2386GAT(755) ,
  \3076GAT(1032)  = ~\3027GAT(1004)  & ~\3026GAT(1003) ,
  \5519GAT(2091)  = ~\5460GAT(2078)  & ~\5459GAT(2065) ,
  \3499GAT(1232)  = ~\3433GAT(1212)  & ~\3377GAT(1189) ,
  \3857GAT(1389)  = ~\3784GAT(1359)  & ~\3628GAT(1289) ,
  \2380GAT(757)  = ~\2339GAT(735)  & ~\2338GAT(730) ,
  \4519GAT(1647)  = ~\4456GAT(1625)  & ~\4398GAT(1596) ,
  \1315GAT(301)  = ~\639GAT(255) ,
  \2265GAT(686)  = ~\2139GAT(625)  & ~\2217GAT(643) ,
  \1594GAT(418)  = ~\1532GAT(392)  & ~\1531GAT(391) ,
  \3458GAT(1202)  = ~\3397GAT(1190)  & ~\3396GAT(1183) ,
  \3764GAT(1364)  = ~\615GAT(263)  & ~\3709GAT(1341) ,
  \1506GAT(406)  = ~\1446GAT(362)  & ~\1401GAT(347) ,
  \5645GAT(2145)  = ~\5575GAT(2119)  & ~\5578GAT(2118) ,
  \2777GAT(917)  = ~\942GAT(154)  & ~\2718GAT(896) ,
  \597GAT(269)  = \307GAT(18)  & \18GAT(1) ,
  \5287GAT(1983)  = ~\5221GAT(1958)  & ~\5160GAT(1934) ,
  \876GAT(176)  = \528GAT(31)  & \103GAT(6) ,
  \6205GAT(2405)  = ~\6201GAT(2402)  & ~\6058GAT(2325) ,
  \5554GAT(2126)  = ~\5489GAT(2109)  & ~\5318GAT(2026) ,
  \1628GAT(439)  = ~\1508GAT(405)  & ~\1582GAT(422) ,
  \5813GAT(2233)  = ~\972GAT(144)  & ~\5761GAT(2199) ,
  \5911GAT(2264)  = ~\5861GAT(2255)  & ~\5810GAT(2222) ,
  \4509GAT(1651)  = ~\4444GAT(1641)  & ~\4281GAT(1555) ,
  \6010GAT(2323)  = ~\5935GAT(2293)  & ~\5975GAT(2307) ,
  \2410GAT(746)  = ~\2359GAT(717)  & ~\1275GAT(43) ,
  \4018GAT(1465)  = ~\3857GAT(1389)  & ~\3971GAT(1437) ,
  \4329GAT(1580)  = ~\4269GAT(1571)  & ~\4085GAT(1479) ,
  \2204GAT(646)  = ~\2129GAT(629)  & ~\2070GAT(610) ,
  \3835GAT(1384)  = ~\3768GAT(1363)  & ~\3712GAT(1339) ,
  \4203GAT(1529)  = ~\4134GAT(1510)  & ~\4070GAT(1483) ,
  \3932GAT(1408)  = ~\3877GAT(1382)  & ~\3693GAT(1299) ,
  \5275GAT(1988)  = ~\5209GAT(1972)  & ~\5148GAT(1937) ,
  \4159GAT(1499)  = ~\4094GAT(1487)  & ~\4040GAT(1446) ,
  \2980GAT(985)  = ~\2922GAT(972)  & ~\2921GAT(966) ,
  \4005GAT(1463)  = ~\3947GAT(1443)  & ~\3896GAT(1422) ,
  \4306GAT(1591)  = ~\4190GAT(1544)  & ~\4251GAT(1566) ,
  \3905GAT(1417)  = ~\3846GAT(1394)  & ~\3845GAT(1381) ,
  \4612GAT(1713)  = ~\4488GAT(1658)  & ~\4557GAT(1679) ,
  \594GAT(270)  = \290GAT(17)  & \18GAT(1) ,
  \2599GAT(857)  = ~\2483GAT(820)  & ~\2552GAT(838) ,
  \2603GAT(856)  = ~\2488GAT(818)  & ~\2555GAT(837) ,
  \3132GAT(1053)  = ~\3016GAT(1007)  & ~\3070GAT(1035) ,
  \4180GAT(1548)  = ~\4114GAT(1515)  & ~\3951GAT(1442) ,
  \4587GAT(1682)  = ~\1251GAT(51)  & ~\4521GAT(1646) ,
  \5993GAT(2301)  = ~\5955GAT(2291)  & ~\5954GAT(2283) ,
  \3026GAT(1003)  = ~\2983GAT(984)  & ~\1281GAT(41) ,
  \4715GAT(1772)  = ~\4541GAT(1694)  & ~\4658GAT(1744) ,
  \1466GAT(357)  = ~\786GAT(206)  & ~\1416GAT(342) ,
  \4634GAT(1704)  = ~\4583GAT(1671)  & ~\4582GAT(1670) ,
  \3398GAT(1182)  = ~\3344GAT(1163)  & ~\3193GAT(1075) ,
  \3336GAT(1169)  = ~\3172GAT(1093)  & ~\3288GAT(1142) ,
  \5840GAT(2257)  = ~\681GAT(241)  & ~\5789GAT(2229) ,
  \5427GAT(2076)  = ~\5370GAT(2057)  & ~\5312GAT(2028) ,
  \2414GAT(782)  = ~\555GAT(283)  & ~\2362GAT(763) ,
  \4167GAT(1496)  = ~\4100GAT(1474)  & ~\4103GAT(1473) ,
  \1343GAT(294)  = ~\975GAT(143) ,
  \5366GAT(2058)  = ~\5241GAT(2008)  & ~\5309GAT(2029) ,
  \1547GAT(383)  = ~\930GAT(158)  & ~\1478GAT(354) ,
  \5249GAT(1995)  = ~\5184GAT(1975)  & ~\5124GAT(1946) ,
  \5984GAT(2311)  = ~\780GAT(208)  & ~\5947GAT(2284) ,
  \3865GAT(1376)  = ~\3793GAT(1357)  & ~\3792GAT(1354) ,
  \4462GAT(1668)  = ~\573GAT(277)  & ~\4405GAT(1643) ,
  \5076GAT(1925)  = ~\819GAT(195)  & ~\5023GAT(1892) ,
  \4575GAT(1673)  = ~\4508GAT(1660)  & ~\4507GAT(1652) ,
  \5954GAT(2283)  = ~\5907GAT(2273)  & ~\5858GAT(2245) ,
  \2996GAT(1027)  = ~\2828GAT(954)  & ~\2942GAT(998) ,
  \3001GAT(1012)  = ~\2954GAT(995)  & ~\2899GAT(975) ,
  \1624GAT(408)  = ~\1578GAT(363)  & ~\1266GAT(46) ,
  \2671GAT(865)  = ~\2631GAT(849)  & ~\2576GAT(830) ,
  \2125GAT(630)  = ~\1032GAT(124)  & ~\2067GAT(612) ,
  \5439GAT(2080)  = ~\822GAT(194)  & ~\5383GAT(2054) ,
  \3847GAT(1393)  = ~\3776GAT(1361)  & ~\3620GAT(1291) ,
  \2905GAT(971)  = ~\2857GAT(938)  & ~\2856GAT(931) ,
  \3883GAT(1370)  = ~\3809GAT(1356)  & ~\3653GAT(1279) ,
  \2942GAT(998)  = ~\2828GAT(954)  & ~\2890GAT(978) ,
  \2273GAT(715)  = ~\2156GAT(680)  & ~\2227GAT(698) ,
  \2264GAT(685)  = ~\2217GAT(643)  & ~\2142GAT(624) ,
  \5063GAT(1879)  = ~\5001GAT(1855)  & ~\1302GAT(34) ,
  \2021GAT(590)  = ~\1866GAT(519)  & ~\1979GAT(569) ,
  \5637GAT(2148)  = ~\5569GAT(2131)  & ~\5507GAT(2094) ,
  \2672GAT(872)  = ~\2523GAT(797)  & ~\2631GAT(849) ,
  \1296GAT(36)  = \460GAT(27)  & \256GAT(15) ,
  \1206GAT(66)  = \494GAT(29)  & \222GAT(13) ,
  \1077GAT(109)  = \307GAT(18)  & \188GAT(11) ,
  \1388GAT(315)  = ~\1343GAT(294) ,
  \4398GAT(1596)  = ~\4349GAT(1584)  & ~\4348GAT(1574) ,
  \6246GAT(2426)  = ~\6237GAT(2419)  & ~\6241GAT(2422) ,
  \4620GAT(1710)  = ~\4566GAT(1689)  & ~\4500GAT(1653) ,
  \2582GAT(827)  = ~\2533GAT(791)  & ~\2536GAT(787) ,
  \2338GAT(730)  = ~\2293GAT(710)  & ~\2242GAT(693) ,
  \4118GAT(1514)  = ~\666GAT(246)  & ~\4058GAT(1489) ,
  \2191GAT(659)  = ~\2117GAT(632)  & ~\1979GAT(569) ,
  \5586GAT(2116)  = ~\5461GAT(2064)  & ~\5522GAT(2090) ,
  \4601GAT(1717)  = ~\4545GAT(1693)  & ~\4544GAT(1683) ,
  \4026GAT(1452)  = ~\3980GAT(1435)  & ~\3923GAT(1410) ,
  \3755GAT(1324)  = ~\3702GAT(1305)  & ~\3659GAT(1276) ,
  \5879GAT(2238)  = ~\5830GAT(2217)  & ~\5829GAT(2216) ,
  \4730GAT(1758)  = ~\4676GAT(1740)  & ~\4675GAT(1735) ,
  \5738GAT(2207)  = ~\5679GAT(2184)  & ~\5621GAT(2153) ,
  \2914GAT(967)  = ~\2869GAT(928)  & ~\2868GAT(927) ,
  \6108GAT(2362)  = ~\6085GAT(2355)  & ~\6005GAT(2324) ,
  \4160GAT(1507)  = ~\1149GAT(85)  & ~\4094GAT(1487) ,
  \1299GAT(35)  = \477GAT(28)  & \256GAT(15) ,
  \1209GAT(65)  = \511GAT(30)  & \222GAT(13) ,
  \4977GAT(1863)  = ~\4921GAT(1843)  & ~\4920GAT(1830) ,
  \4947GAT(1875)  = ~\4885GAT(1852)  & ~\4884GAT(1841) ,
  \5522GAT(2090)  = ~\5461GAT(2064)  & ~\5464GAT(2063) ,
  \624GAT(260)  = \460GAT(27)  & \18GAT(1) ,
  \5526GAT(2088)  = ~\5467GAT(2062)  & ~\5413GAT(2039) ,
  \6157GAT(2379)  = ~\6151GAT(2377)  & ~\6114GAT(2359) ,
  \2186GAT(662)  = ~\2113GAT(633)  & ~\1975GAT(570) ,
  \4896GAT(1847)  = ~\4829GAT(1818)  & ~\4658GAT(1744) ,
  \4435GAT(1632)  = ~\4374GAT(1604)  & ~\4377GAT(1603) ,
  \1546GAT(382)  = ~\1478GAT(354)  & ~\1425GAT(339) ,
  \2781GAT(916)  = ~\990GAT(138)  & ~\2721GAT(895) ,
  \5115GAT(1903)  = ~\5064GAT(1880)  & ~\5063GAT(1879) ,
  \2492GAT(817)  = ~\699GAT(235)  & ~\2426GAT(779) ,
  \2190GAT(661)  = ~\936GAT(156)  & ~\2117GAT(632) ,
  \5501GAT(2097)  = ~\5440GAT(2071)  & ~\5443GAT(2070) ,
  \1290GAT(38)  = \426GAT(25)  & \256GAT(15) ,
  \1293GAT(37)  = \443GAT(26)  & \256GAT(15) ,
  \1203GAT(67)  = \477GAT(28)  & \222GAT(13) ,
  \1200GAT(68)  = \460GAT(27)  & \222GAT(13) ,
  \5378GAT(2050)  = ~\5318GAT(2026)  & ~\5259GAT(1993) ,
  \5782GAT(2192)  = ~\5726GAT(2169)  & ~\5725GAT(2168) ,
  \4079GAT(1481)  = ~\4022GAT(1464)  & ~\3868GAT(1375) ,
  \546GAT(286)  = \290GAT(17)  & \1GAT(0) ,
  \6073GAT(2341)  = ~\6045GAT(2334)  & ~\6044GAT(2331) ,
  \6147GAT(2374)  = ~\6141GAT(2373)  & ~\6124GAT(2367) ,
  \2511GAT(795)  = ~\2442GAT(775)  & ~\2383GAT(756) ,
  \930GAT(158)  = \290GAT(17)  & \137GAT(8) ,
  \4838GAT(1816)  = ~\816GAT(196)  & ~\4775GAT(1798) ,
  \1437GAT(335)  = ~\1396GAT(307)  & ~\1395GAT(308) ,
  \2950GAT(996)  = ~\2838GAT(948)  & ~\2896GAT(976) ,
  \4531GAT(1698)  = ~\4466GAT(1667)  & ~\4298GAT(1593) ,
  \2242GAT(693)  = ~\2185GAT(664)  & ~\2184GAT(657) ,
  \3480GAT(1254)  = ~\564GAT(280)  & ~\3417GAT(1216) ,
  \1389GAT(314)  = ~\1347GAT(293)  & ~\1023GAT(127) ,
  \2917GAT(974)  = ~\1185GAT(73)  & ~\2870GAT(926) ,
  \4886GAT(1851)  = ~\4821GAT(1820)  & ~\4650GAT(1746) ,
  \1756GAT(469)  = ~\1713GAT(442)  & ~\1712GAT(441) ,
  \1351GAT(292)  = ~\1071GAT(111) ,
  \2383GAT(756)  = ~\2341GAT(733)  & ~\2340GAT(728) ,
  \2649GAT(845)  = ~\1230GAT(58)  & ~\2591GAT(829) ,
  \2724GAT(894)  = ~\2674GAT(870)  & ~\2673GAT(864) ,
  \2339GAT(735)  = ~\2181GAT(665)  & ~\2293GAT(710) ,
  \1434GAT(336)  = ~\1394GAT(309)  & ~\1393GAT(310) ,
  \1597GAT(417)  = ~\1537GAT(389)  & ~\1536GAT(388) ,
  \2085GAT(640)  = ~\552GAT(284)  & ~\2037GAT(622) ,
  \4189GAT(1545)  = ~\714GAT(230)  & ~\4122GAT(1513) ,
  \3453GAT(1204)  = ~\3392GAT(1192)  & ~\3341GAT(1156) ,
  \768GAT(212)  = \460GAT(27)  & \69GAT(4) ,
  \4985GAT(1861)  = ~\4860GAT(1804)  & ~\4928GAT(1827) ,
  \5870GAT(2242)  = ~\5818GAT(2232)  & ~\5817GAT(2221) ,
  \5611GAT(2155)  = ~\5544GAT(2134)  & ~\5483GAT(2103) ,
  \1011GAT(131)  = \477GAT(28)  & \154GAT(9) ,
  \4683GAT(1732)  = ~\4622GAT(1709)  & ~\4625GAT(1708) ,
  \1791GAT(493)  = ~\885GAT(173)  & ~\1738GAT(476) ,
  \4174GAT(1551)  = ~\570GAT(278)  & ~\4110GAT(1516) ,
  \5262GAT(1992)  = ~\5194GAT(1967)  & ~\5197GAT(1966) ,
  \3501GAT(1245)  = ~\3433GAT(1212)  & ~\3280GAT(1144) ,
  \630GAT(258)  = \494GAT(29)  & \18GAT(1) ,
  \4708GAT(1768)  = ~\4646GAT(1747)  & ~\4592GAT(1721) ,
  \561GAT(281)  = \375GAT(22)  & \1GAT(0) ,
  \1390GAT(313)  = ~\1347GAT(293) ,
  \5856GAT(2246)  = ~\5804GAT(2225)  & ~\5752GAT(2203) ,
  \849GAT(185)  = \375GAT(22)  & \103GAT(6) ,
  \5147GAT(1939)  = ~\5032GAT(1890)  & ~\5088GAT(1913) ,
  \545GAT(287)  = \[0] ,
  \5288GAT(1984)  = ~\5157GAT(1935)  & ~\5221GAT(1958) ,
  \1963GAT(573)  = ~\1846GAT(531)  & ~\1914GAT(556) ,
  \2670GAT(874)  = ~\2518GAT(800)  & ~\2627GAT(850) ,
  \2673GAT(864)  = ~\2635GAT(848)  & ~\2579GAT(828) ,
  \4907GAT(1834)  = ~\4839GAT(1811)  & ~\4842GAT(1810) ,
  \5080GAT(1916)  = ~\5026GAT(1897)  & ~\4965GAT(1866) ,
  \6045GAT(2334)  = ~\732GAT(224)  & ~\6014GAT(2322) ,
  \627GAT(259)  = \477GAT(28)  & \18GAT(1) ,
  \1044GAT(120)  = \392GAT(23)  & \171GAT(10) ,
  \2350GAT(719)  = ~\2318GAT(704)  & ~\2317GAT(702) ,
  \2113GAT(633)  = ~\888GAT(172)  & ~\2058GAT(615) ,
  \3571GAT(1266)  = ~\3515GAT(1239)  & ~\3514GAT(1227) ,
  \6221GAT(2412)  = ~\6217GAT(2409)  & ~\6002GAT(2297) ,
  \1281GAT(41)  = \375GAT(22)  & \256GAT(15) ,
  \1221GAT(61)  = \307GAT(18)  & \239GAT(14) ,
  \3583GAT(1261)  = ~\3532GAT(1223)  & ~\3531GAT(1222) ,
  \2475GAT(765)  = ~\2359GAT(717)  & ~\2410GAT(746) ,
  \2493GAT(815)  = ~\2426GAT(779)  & ~\2281GAT(713) ,
  \1319GAT(300)  = ~\687GAT(239) ,
  \5430GAT(2082)  = ~\5251GAT(2004)  & ~\5374GAT(2056) ,
  \2023GAT(588)  = ~\1871GAT(516)  & ~\1983GAT(568) ,
  \2816GAT(949)  = ~\2753GAT(923)  & ~\2700GAT(904) ,
  \2861GAT(930)  = ~\2790GAT(914)  & ~\2789GAT(913) ,
  \2648GAT(842)  = ~\2591GAT(829)  & ~\2545GAT(783) ,
  \2189GAT(654)  = ~\2117GAT(632)  & ~\2061GAT(614) ,
  \1284GAT(40)  = \392GAT(23)  & \256GAT(15) ,
  \1224GAT(60)  = \324GAT(19)  & \239GAT(14) ,
  \3349GAT(1161)  = ~\1092GAT(104)  & ~\3305GAT(1138) ,
  \5255GAT(2003)  = ~\723GAT(227)  & ~\5188GAT(1974) ,
  \3309GAT(1134)  = ~\3248GAT(1121)  & ~\3199GAT(1072) ,
  \2336GAT(732)  = ~\2289GAT(711)  & ~\2239GAT(694) ,
  \4739GAT(1754)  = ~\4688GAT(1731)  & ~\4687GAT(1730) ,
  \3146GAT(1106)  = ~\609GAT(265)  & ~\3083GAT(1068) ,
  \4760GAT(1795)  = ~\4709GAT(1775)  & ~\4708GAT(1768) ,
  \2555GAT(837)  = ~\2492GAT(817)  & ~\2491GAT(807) ,
  \4875GAT(1813)  = ~\1254GAT(50)  & ~\4814GAT(1776) ,
  \1391GAT(312)  = ~\1351GAT(292)  & ~\1071GAT(111) ,
  \2337GAT(737)  = ~\2176GAT(668)  & ~\2289GAT(711) ,
  \2908GAT(970)  = ~\2858GAT(936)  & ~\2861GAT(930) ,
  \1287GAT(39)  = \409GAT(24)  & \256GAT(15) ,
  \1272GAT(44)  = \324GAT(19)  & \256GAT(15) ,
  \1227GAT(59)  = \341GAT(20)  & \239GAT(14) ,
  \1212GAT(64)  = \528GAT(31)  & \222GAT(13) ,
  \5483GAT(2103)  = ~\5428GAT(2083)  & ~\5427GAT(2076) ,
  \5837GAT(2252)  = ~\5788GAT(2236)  & ~\5787GAT(2230) ,
  \5996GAT(2300)  = ~\5956GAT(2282)  & ~\5959GAT(2281) ,
  \3697GAT(1297)  = ~\3653GAT(1279)  & ~\3595GAT(1258) ,
  \717GAT(229)  = \443GAT(26)  & \52GAT(3) ,
  \6119GAT(2358)  = ~\6070GAT(2342)  & ~\6097GAT(2350) ,
  \2666GAT(878)  = ~\2508GAT(806)  & ~\2619GAT(852) ,
  \2418GAT(781)  = ~\603GAT(267)  & ~\2365GAT(762) ,
  \5845GAT(2256)  = ~\729GAT(225)  & ~\5792GAT(2235) ,
  \5476GAT(2075)  = ~\1260GAT(48)  & ~\5422GAT(2035) ,
  \969GAT(145)  = \511GAT(30)  & \137GAT(8) ,
  \6135GAT(2369)  = ~\6129GAT(2366)  & ~\6128GAT(2365) ,
  \5395GAT(2045)  = ~\5333GAT(2021)  & ~\5336GAT(2020) ,
  \4837GAT(1812)  = ~\4775GAT(1798)  & ~\4718GAT(1761) ,
  \1581GAT(423)  = \[1] ,
  \3162GAT(1099)  = ~\3095GAT(1065)  & ~\2942GAT(998) ,
  \2790GAT(914)  = ~\1086GAT(106)  & ~\2727GAT(899) ,
  \1392GAT(311)  = ~\1351GAT(292) ,
  \1384GAT(319)  = ~\1335GAT(296) ,
  \4641GAT(1703)  = ~\4587GAT(1682)  & ~\4521GAT(1646) ,
  \2474GAT(764)  = ~\2410GAT(746)  & ~\1275GAT(43) ,
  \2811GAT(952)  = ~\2749GAT(924)  & ~\2697GAT(905) ,
  \4070GAT(1483)  = ~\4018GAT(1465)  & ~\4017GAT(1454) ,
  \1278GAT(42)  = \358GAT(21)  & \256GAT(15) ,
  \1218GAT(62)  = \290GAT(17)  & \239GAT(14) ,
  \2070GAT(610)  = ~\2027GAT(584)  & ~\2026GAT(581) ,
  \2481GAT(813)  = ~\2418GAT(781)  & ~\2365GAT(762) ,
  \3516GAT(1237)  = ~\3445GAT(1209)  & ~\3292GAT(1141) ,
  \3417GAT(1216)  = ~\564GAT(280)  & ~\3365GAT(1195) ,
  \1047GAT(119)  = \409GAT(24)  & \171GAT(10) ,
  \2727GAT(899)  = ~\1086GAT(106)  & ~\2675GAT(863) ,
  \4287GAT(1552)  = ~\4237GAT(1519)  & ~\4236GAT(1518) ,
  \714GAT(230)  = \426GAT(25)  & \52GAT(3) ,
  \3330GAT(1173)  = ~\3157GAT(1101)  & ~\3276GAT(1145) ,
  \4633GAT(1706)  = ~\4509GAT(1651)  & ~\4578GAT(1672) ,
  \1275GAT(43)  = \341GAT(20)  & \256GAT(15) ,
  \1215GAT(63)  = \273GAT(16)  & \239GAT(14) ,
  \4275GAT(1557)  = ~\4220GAT(1535)  & ~\4034GAT(1449) ,
  \5452GAT(2066)  = ~\5400GAT(2044)  & ~\5399GAT(2043) ,
  \4393GAT(1598)  = ~\4344GAT(1585)  & ~\4287GAT(1552) ,
  \4245GAT(1568)  = ~\4184GAT(1547)  & ~\4183GAT(1534) ,
  \4363GAT(1607)  = ~\4314GAT(1589)  & ~\4257GAT(1563) ,
  \3397GAT(1190)  = ~\1044GAT(120)  & ~\3344GAT(1163) ,
  \1741GAT(475)  = ~\1703GAT(452)  & ~\1702GAT(451) ,
  \4849GAT(1807)  = ~\4787GAT(1786)  & ~\4730GAT(1758) ,
  \4525GAT(1701)  = ~\573GAT(277)  & ~\4462GAT(1668) ,
  \2813GAT(961)  = ~\2749GAT(924)  & ~\2599GAT(857) ,
  \933GAT(157)  = \307GAT(18)  & \137GAT(8) ,
  \5704GAT(2175)  = ~\5645GAT(2145)  & ~\5578GAT(2118) ,
  \5259GAT(1993)  = ~\5193GAT(1973)  & ~\5192GAT(1968) ,
  \4205GAT(1538)  = ~\4134GAT(1510)  & ~\3971GAT(1437) ,
  \4385GAT(1601)  = ~\4275GAT(1557)  & ~\4335GAT(1578) ,
  \1266GAT(46)  = \290GAT(17)  & \256GAT(15) ,
  \1236GAT(56)  = \392GAT(23)  & \239GAT(14) ,
  \4038GAT(1447)  = ~\3992GAT(1427)  & ~\3935GAT(1407) ,
  \3107GAT(1062)  = ~\897GAT(169)  & ~\3049GAT(1041) ,
  \2483GAT(820)  = ~\2418GAT(781)  & ~\2273GAT(715) ,
  \2022GAT(585)  = ~\1983GAT(568)  & ~\1929GAT(551) ,
  \5051GAT(1884)  = ~\4989GAT(1874)  & ~\4934GAT(1824) ,
  \5566GAT(2121)  = ~\5506GAT(2096)  & ~\5505GAT(2095) ,
  \4224GAT(1523)  = ~\4155GAT(1508)  & ~\4091GAT(1476) ,
  \5245GAT(2007)  = ~\627GAT(259)  & ~\5180GAT(1976) ,
  \3239GAT(1116)  = ~\3187GAT(1084)  & ~\3190GAT(1076) ,
  \1393GAT(310)  = ~\1355GAT(291)  & ~\1119GAT(95) ,
  \1385GAT(318)  = ~\1339GAT(295)  & ~\927GAT(159) ,
  \2791GAT(912)  = ~\2727GAT(899)  & ~\2582GAT(827) ,
  \6076GAT(2340)  = ~\6046GAT(2330)  & ~\6049GAT(2329) ,
  \2334GAT(734)  = ~\2285GAT(712)  & ~\2236GAT(695) ,
  \5537GAT(2085)  = ~\5476GAT(2075)  & ~\5304GAT(1978) ,
  \4139GAT(1509)  = ~\906GAT(166)  & ~\4073GAT(1493) ,
  \3485GAT(1252)  = ~\612GAT(264)  & ~\3421GAT(1215) ,
  \1269GAT(45)  = \307GAT(18)  & \256GAT(15) ,
  \1239GAT(55)  = \409GAT(24)  & \239GAT(14) ,
  \3495GAT(1248)  = ~\708GAT(232)  & ~\3429GAT(1213) ,
  \5788GAT(2236)  = ~\5613GAT(2163)  & ~\5734GAT(2213) ,
  \3959GAT(1440)  = ~\3842GAT(1395)  & ~\3905GAT(1417) ,
  \3140GAT(1097)  = ~\3079GAT(1069)  & ~\3028GAT(1050) ,
  \5148GAT(1937)  = ~\5093GAT(1912)  & ~\5092GAT(1911) ,
  \1074GAT(110)  = \290GAT(17)  & \188GAT(11) ,
  \1911GAT(557)  = ~\1845GAT(533)  & ~\1844GAT(529) ,
  \2335GAT(739)  = ~\2171GAT(671)  & ~\2285GAT(712) ,
  \5715GAT(2172)  = ~\5654GAT(2158)  & ~\5467GAT(2062) ,
  \4710GAT(1766)  = ~\4650GAT(1746)  & ~\4595GAT(1720) ,
  \633GAT(257)  = \511GAT(30)  & \18GAT(1) ,
  \2491GAT(807)  = ~\2426GAT(779)  & ~\2371GAT(760) ,
  \3914GAT(1414)  = ~\3861GAT(1388)  & ~\3860GAT(1377) ,
  \3064GAT(1037)  = ~\3010GAT(1015)  & ~\2864GAT(929) ,
  \1263GAT(47)  = \273GAT(16)  & \256GAT(15) ,
  \1260GAT(48)  = \528GAT(31)  & \239GAT(14) ,
  \1233GAT(57)  = \375GAT(22)  & \239GAT(14) ,
  \1230GAT(58)  = \358GAT(21)  & \239GAT(14) ,
  \3886GAT(1369)  = ~\3814GAT(1355)  & ~\3813GAT(1347) ,
  \4688GAT(1731)  = ~\4572GAT(1674)  & ~\4628GAT(1707) ,
  \6165GAT(2385)  = ~\6161GAT(2382)  & ~\6130GAT(2364) ,
  \1709GAT(446)  = ~\1563GAT(372)  & ~\1672GAT(428) ,
  \5109GAT(1906)  = ~\5053GAT(1883)  & ~\5056GAT(1882) ,
  \3034GAT(1048)  = ~\2992GAT(1029)  & ~\2991GAT(1022) ,
  \1257GAT(49)  = \511GAT(30)  & \239GAT(14) ,
  \1242GAT(54)  = \426GAT(25)  & \239GAT(14) ,
  \2353GAT(723)  = ~\1179GAT(75)  & ~\2319GAT(701) ,
  \1508GAT(405)  = ~\1446GAT(362)  & ~\1311GAT(302) ,
  \5312GAT(2028)  = ~\5250GAT(2005)  & ~\5249GAT(1995) ,
  \4354GAT(1622)  = ~\4175GAT(1550)  & ~\4294GAT(1594) ,
  \1577GAT(365)  = ~\1218GAT(62)  & ~\1502GAT(348) ,
  \2667GAT(869)  = ~\2623GAT(851)  & ~\2570GAT(832) ,
  \2482GAT(821)  = ~\603GAT(267)  & ~\2418GAT(781) ,
  \4440GAT(1631)  = ~\4329GAT(1580)  & ~\4380GAT(1602) ,
  \3206GAT(1071)  = ~\3136GAT(1058)  & ~\3076GAT(1032) ,
  \3568GAT(1267)  = ~\3510GAT(1242)  & ~\3509GAT(1229) ,
  \3360GAT(1150)  = ~\3317GAT(1131)  & ~\3257GAT(1110) ,
  \1443GAT(333)  = ~\1400GAT(303)  & ~\1399GAT(304) ,
  \5902GAT(2266)  = ~\5852GAT(2248)  & ~\5801GAT(2226) ,
  \2301GAT(708)  = ~\2191GAT(659)  & ~\2248GAT(691) ,
  \3659GAT(1276)  = ~\3603GAT(1256)  & ~\3602GAT(1255) ,
  \5283GAT(1985)  = ~\5215GAT(1960)  & ~\5218GAT(1959) ,
  \3467GAT(1198)  = ~\3409GAT(1179)  & ~\3408GAT(1178) ,
  \6120GAT(2356)  = ~\6102GAT(2349)  & ~\6101GAT(2348) ,
  \2812GAT(962)  = ~\606GAT(266)  & ~\2749GAT(924) ,
  \4860GAT(1804)  = ~\4796GAT(1796)  & ~\4628GAT(1707) ,
  \4091GAT(1476)  = ~\4039GAT(1448)  & ~\4038GAT(1447) ,
  \1248GAT(52)  = \460GAT(27)  & \239GAT(14) ,
  \6270GAT(2438)  = \[28] ,
  \1386GAT(317)  = ~\1339GAT(295) ,
  \5127GAT(1944)  = ~\5072GAT(1926)  & ~\5071GAT(1918) ,
  \5157GAT(1935)  = ~\5097GAT(1923)  & ~\4928GAT(1827) ,
  \5510GAT(2107)  = ~\969GAT(145)  & ~\5452GAT(2066) ,
  \3302GAT(1135)  = ~\3244GAT(1115)  & ~\3243GAT(1114) ,
  \2020GAT(587)  = ~\1979GAT(569)  & ~\1926GAT(552) ,
  \741GAT(221)  = \307GAT(18)  & \69GAT(4) ,
  \1339GAT(295)  = ~\927GAT(159) ,
  \3645GAT(1282)  = ~\3586GAT(1270)  & ~\3533GAT(1221) ,
  \966GAT(146)  = \494GAT(29)  & \137GAT(8) ,
  \3454GAT(1207)  = ~\996GAT(136)  & ~\3392GAT(1192) ,
  \1562GAT(374)  = ~\1074GAT(110)  & ~\1490GAT(351) ,
  \2463GAT(770)  = ~\1131GAT(91)  & ~\2398GAT(754) ,
  \5336GAT(2020)  = ~\5276GAT(2000)  & ~\5275GAT(1988) ,
  \1245GAT(53)  = \443GAT(26)  & \239GAT(14) ,
  \5849GAT(2249)  = ~\5797GAT(2234)  & ~\5796GAT(2228) ,
  \4607GAT(1714)  = ~\4551GAT(1690)  & ~\4554GAT(1680) ,
  \1759GAT(470)  = ~\1221GAT(61)  & ~\1714GAT(440) ,
  \2644GAT(846)  = ~\1182GAT(74)  & ~\2588GAT(824) ,
  \3466GAT(1200)  = ~\3350GAT(1154)  & ~\3404GAT(1180) ,
  \4769GAT(1791)  = ~\4715GAT(1772)  & ~\4714GAT(1763) ,
  \4792GAT(1785)  = ~\4677GAT(1734)  & ~\4733GAT(1757) ,
  \5197GAT(1966)  = ~\5135GAT(1951)  & ~\5134GAT(1943) ,
  \3010GAT(1015)  = ~\1089GAT(105)  & ~\2968GAT(988) ,
  \4014GAT(1467)  = ~\3847GAT(1393)  & ~\3963GAT(1439) ,
  \3746GAT(1326)  = ~\3693GAT(1299)  & ~\3650GAT(1280) ,
  \1008GAT(132)  = \460GAT(27)  & \154GAT(9) ,
  \3063GAT(1043)  = ~\1089GAT(105)  & ~\3010GAT(1015) ,
  \4200GAT(1540)  = ~\4130GAT(1511)  & ~\3967GAT(1438) ,
  \555GAT(283)  = \341GAT(20)  & \1GAT(0) ,
  \1176GAT(76)  = \324GAT(19)  & \222GAT(13) ,
  \1440GAT(334)  = ~\1398GAT(305)  & ~\1397GAT(306) ,
  \3120GAT(1059)  = ~\1041GAT(121)  & ~\3058GAT(1045) ,
  \1576GAT(364)  = ~\1502GAT(348)  & ~\1443GAT(333) ,
  \687GAT(239)  = \273GAT(16)  & \52GAT(3) ,
  \4152GAT(1500)  = ~\4090GAT(1478)  & ~\4089GAT(1477) ,
  \819GAT(195)  = \477GAT(28)  & \86GAT(5) ,
  \1582GAT(422)  = ~\1512GAT(404)  & ~\1511GAT(403) ,
  \5308GAT(2031)  = \[12] ,
  \1548GAT(381)  = ~\1478GAT(354)  & ~\1343GAT(294) ,
  \879GAT(175)  = \273GAT(16)  & \120GAT(7) ,
  \2721GAT(895)  = ~\2672GAT(872)  & ~\2671GAT(865) ,
  \3014GAT(1008)  = ~\2971GAT(991)  & ~\2914GAT(967) ,
  \3826GAT(1402)  = ~\567GAT(279)  & ~\3760GAT(1365) ,
  \5206GAT(1962)  = ~\5147GAT(1939)  & ~\5146GAT(1938) ,
  \4879GAT(1842)  = ~\4817GAT(1821)  & ~\4760GAT(1795) ,
  \3975GAT(1432)  = ~\3917GAT(1413)  & ~\3865GAT(1376) ,
  \4704GAT(1725)  = ~\4643GAT(1702)  & ~\1299GAT(35) ,
  \4994GAT(1872)  = ~\1206GAT(66)  & ~\4937GAT(1839) ,
  \1502GAT(348)  = ~\1218GAT(62)  & ~\1443GAT(333) ,
  \549GAT(285)  = \307GAT(18)  & \1GAT(0) ,
  \5923GAT(2259)  = ~\5873GAT(2241)  & ~\5822GAT(2219) ,
  \3156GAT(1102)  = ~\705GAT(233)  & ~\3091GAT(1066) ,
  \1708GAT(445)  = ~\1672GAT(428)  & ~\1615GAT(411) ,
  \765GAT(213)  = \443GAT(26)  & \69GAT(4) ,
  \6185GAT(2395)  = ~\6181GAT(2392)  & ~\6103GAT(2347) ,
  \1387GAT(316)  = ~\1343GAT(294)  & ~\975GAT(143) ,
  \1179GAT(75)  = \341GAT(20)  & \222GAT(13) ,
  \4549GAT(1681)  = ~\4482GAT(1663)  & ~\4420GAT(1636) ,
  \2665GAT(871)  = ~\2619GAT(852)  & ~\2567GAT(833) ,
  \6226GAT(2416)  = ~\6217GAT(2409)  & ~\6221GAT(2412) ,
  \4067GAT(1484)  = ~\4016GAT(1466)  & ~\4015GAT(1456) ,
  \6171GAT(2387)  = ~\6167GAT(2384)  & ~\6120GAT(2356) ,
  \1874GAT(511)  = ~\1803GAT(490)  & ~\1747GAT(473) ,
  \2664GAT(880)  = ~\2503GAT(809)  & ~\2615GAT(853) ,
  \3967GAT(1438)  = ~\3852GAT(1391)  & ~\3911GAT(1415) ,
  \3793GAT(1357)  = ~\951GAT(151)  & ~\3730GAT(1342) ,
  \5505GAT(2095)  = ~\5446GAT(2069)  & ~\5392GAT(2046) ,
  \3005GAT(1010)  = ~\2962GAT(993)  & ~\2905GAT(971) ,
  \4545GAT(1693)  = ~\765GAT(213)  & ~\4478GAT(1664) ,
  \6287GAT(2444)  = \[30] ,
  \3542GAT(1219)  = ~\3470GAT(1206)  & ~\3317GAT(1131) ,
  \4427GAT(1635)  = ~\4368GAT(1616)  & ~\4320GAT(1582) ,
  \945GAT(153)  = \375GAT(22)  & \137GAT(8) ,
  \2340GAT(728)  = ~\2297GAT(709)  & ~\2245GAT(692) ,
  \3136GAT(1058)  = ~\1236GAT(56)  & ~\3076GAT(1032) ,
  \1707GAT(448)  = ~\1558GAT(375)  & ~\1668GAT(429) ,
  \4236GAT(1518)  = ~\4167GAT(1496)  & ~\4103GAT(1473) ,
  \1563GAT(372)  = ~\1490GAT(351)  & ~\1355GAT(291) ,
  \1173GAT(77)  = \307GAT(18)  & \222GAT(13) ,
  \1170GAT(78)  = \290GAT(17)  & \222GAT(13) ,
  \4671GAT(1741)  = ~\912GAT(164)  & ~\4613GAT(1711) ,
  \4989GAT(1874)  = ~\1158GAT(82)  & ~\4934GAT(1824) ,
  \3181GAT(1089)  = ~\945GAT(153)  & ~\3111GAT(1061) ,
  \5486GAT(2101)  = ~\5430GAT(2082)  & ~\5429GAT(2074) ,
  \5907GAT(2273)  = ~\876GAT(176)  & ~\5858GAT(2245) ,
  \3650GAT(1280)  = ~\3591GAT(1268)  & ~\3590GAT(1260) ,
  \2588GAT(824)  = ~\2544GAT(785)  & ~\2543GAT(784) ,
  \1182GAT(74)  = \358GAT(21)  & \222GAT(13) ,
  \5072GAT(1926)  = ~\4896GAT(1847)  & ~\5017GAT(1899) ,
  \2073GAT(608)  = ~\2029GAT(582)  & ~\2028GAT(579) ,
  \5928GAT(2290)  = ~\5882GAT(2276)  & ~\5834GAT(2253) ,
  \5890GAT(2271)  = ~\5840GAT(2257)  & ~\5789GAT(2229) ,
  \2869GAT(928)  = ~\2733GAT(892)  & ~\2797GAT(910) ,
  \4916GAT(1844)  = ~\963GAT(147)  & ~\4851GAT(1806) ,
  \2462GAT(769)  = ~\2398GAT(754)  & ~\2350GAT(719) ,
  \4781GAT(1788)  = ~\4721GAT(1770)  & ~\4557GAT(1679) ,
  \843GAT(187)  = \341GAT(20)  & \103GAT(6) ,
  \5498GAT(2098)  = ~\5439GAT(2080)  & ~\5438GAT(2072) ,
  \2343GAT(731)  = ~\2191GAT(659)  & ~\2301GAT(708) ,
  \1446GAT(362)  = ~\546GAT(286)  & ~\1401GAT(347) ,
  \4341GAT(1575)  = ~\4286GAT(1554)  & ~\4285GAT(1553) ,
  \2669GAT(867)  = ~\2627GAT(850)  & ~\2573GAT(831) ,
  \3296GAT(1140)  = ~\3182GAT(1087)  & ~\3236GAT(1117) ,
  \5514GAT(2093)  = ~\5455GAT(2079)  & ~\5401GAT(2042) ,
  \1735GAT(477)  = ~\1699GAT(456)  & ~\1698GAT(455) ,
  \4294GAT(1594)  = ~\4175GAT(1550)  & ~\4242GAT(1570) ,
  \4965GAT(1866)  = ~\4912GAT(1833)  & ~\4911GAT(1832) ,
  \1676GAT(427)  = ~\1568GAT(369)  & ~\1618GAT(410) ,
  \1188GAT(72)  = \392GAT(23)  & \222GAT(13) ,
  \3321GAT(1129)  = ~\3260GAT(1109)  & ~\1284GAT(40) ,
  \3519GAT(1226)  = ~\3449GAT(1208)  & ~\3389GAT(1184) ,
  \6275GAT(2440)  = ~\6271GAT(2437)  & ~\5782GAT(2192) ,
  \1474GAT(355)  = ~\882GAT(174)  & ~\1422GAT(340) ,
  \2498GAT(812)  = ~\2430GAT(778)  & ~\2285GAT(712) ,
  \1975GAT(570)  = ~\1861GAT(522)  & ~\1923GAT(553) ,
  \4941GAT(1823)  = ~\4875GAT(1813)  & ~\4814GAT(1776) ,
  \1700GAT(453)  = ~\1656GAT(432)  & ~\1603GAT(415) ,
  \3996GAT(1425)  = ~\3938GAT(1406)  & ~\3886GAT(1369) ,
  \4439GAT(1630)  = ~\4380GAT(1602)  & ~\4332GAT(1579) ,
  \5792GAT(2235)  = ~\729GAT(225)  & ~\5740GAT(2206) ,
  \5966GAT(2278)  = ~\5919GAT(2261)  & ~\5870GAT(2242) ,
  \4842GAT(1810)  = ~\4780GAT(1797)  & ~\4779GAT(1789) ,
  \6133GAT(2370)  = ~\6124GAT(2367)  & ~\6111GAT(2360) ,
  \1612GAT(412)  = ~\1562GAT(374)  & ~\1561GAT(373) ,
  \2821GAT(946)  = ~\2757GAT(922)  & ~\2703GAT(903) ,
  \1185GAT(73)  = \375GAT(22)  & \222GAT(13) ,
  \3510GAT(1242)  = ~\852GAT(184)  & ~\3441GAT(1210) ,
  \4488GAT(1658)  = ~\4423GAT(1645)  & ~\4260GAT(1562) ,
  \3329GAT(1164)  = ~\3276GAT(1145)  & ~\3221GAT(1124) ,
  \[10]  = ~\4525GAT(1701)  & ~\4524GAT(1688) ,
  \1706GAT(447)  = ~\1668GAT(429)  & ~\1612GAT(412) ,
  \4933GAT(1826)  = ~\4802GAT(1781)  & ~\4866GAT(1802) ,
  \[11]  = ~\4880GAT(1854)  & ~\4879GAT(1842) ,
  \1875GAT(515)  = ~\1029GAT(125)  & ~\1803GAT(490) ,
  \792GAT(204)  = \324GAT(19)  & \86GAT(5) ,
  \4817GAT(1821)  = ~\576GAT(276)  & ~\4760GAT(1795) ,
  \[12]  = ~\5240GAT(2009)  & ~\5239GAT(1999) ,
  \2040GAT(621)  = ~\2007GAT(604)  & ~\2006GAT(601) ,
  \5268GAT(1989)  = ~\5205GAT(1964)  & ~\5204GAT(1963) ,
  \2528GAT(794)  = ~\2454GAT(772)  & ~\2309GAT(706) ,
  \[13]  = ~\5607GAT(2166)  & ~\5606GAT(2156) ,
  \1979GAT(569)  = ~\1866GAT(519)  & ~\1926GAT(552) ,
  \4008GAT(1470)  = ~\3832GAT(1399)  & ~\3951GAT(1442) ,
  \[14]  = ~\5929GAT(2296)  & ~\5928GAT(2290) ,
  \2239GAT(694)  = ~\2180GAT(667)  & ~\2179GAT(660) ,
  \4130GAT(1511)  = ~\810GAT(198)  & ~\4067GAT(1484) ,
  \2868GAT(927)  = ~\2797GAT(910)  & ~\2736GAT(891) ,
  \[15]  = ~\6107GAT(2363)  & ~\6106GAT(2361) ,
  \3489GAT(1235)  = ~\3425GAT(1214)  & ~\3371GAT(1193) ,
  \2526GAT(789)  = ~\2454GAT(772)  & ~\2392GAT(751) ,
  \[16]  = ~\6146GAT(2376)  & ~\6145GAT(2375) ,
  \1879GAT(508)  = ~\1807GAT(489)  & ~\1750GAT(472) ,
  \1578GAT(363)  = ~\1502GAT(348)  & ~\1367GAT(288) ,
  \[17]  = ~\6156GAT(2381)  & ~\6155GAT(2380) ,
  \4314GAT(1589)  = ~\4200GAT(1540)  & ~\4257GAT(1563) ,
  \5225GAT(1956)  = ~\5163GAT(1933)  & ~\5106GAT(1907) ,
  \3943GAT(1405)  = ~\3815GAT(1346)  & ~\3889GAT(1368) ,
  \[18]  = ~\6166GAT(2386)  & ~\6165GAT(2385) ,
  \1161GAT(81)  = \511GAT(30)  & \205GAT(12) ,
  \6081GAT(2339)  = ~\6020GAT(2317)  & ~\6052GAT(2328) ,
  \[19]  = ~\6176GAT(2391)  & ~\6175GAT(2390) ,
  \2496GAT(804)  = ~\2430GAT(778)  & ~\2374GAT(759) ,
  \1701GAT(454)  = ~\1543GAT(384)  & ~\1656GAT(432) ,
  \807GAT(199)  = \409GAT(24)  & \86GAT(5) ,
  \5924GAT(2260)  = ~\5819GAT(2220)  & ~\5873GAT(2241) ,
  \1164GAT(80)  = \528GAT(31)  & \205GAT(12) ,
  \2991GAT(1022)  = ~\2934GAT(1000)  & ~\2884GAT(980) ,
  \4766GAT(1792)  = ~\4713GAT(1773)  & ~\4712GAT(1764) ,
  \2631GAT(849)  = ~\2523GAT(797)  & ~\2576GAT(830) ,
  \750GAT(218)  = \358GAT(21)  & \69GAT(4) ,
  \3756GAT(1333)  = ~\1242GAT(54)  & ~\3702GAT(1305) ,
  \2827GAT(956)  = ~\750GAT(218)  & ~\2761GAT(921) ,
  \5916GAT(2262)  = ~\5866GAT(2254)  & ~\5865GAT(2244) ,
  \684GAT(240)  = \528GAT(31)  & \35GAT(2) ,
  \3150GAT(1091)  = ~\3087GAT(1067)  & ~\3034GAT(1048) ,
  \1561GAT(373)  = ~\1490GAT(351)  & ~\1434GAT(336) ,
  \3908GAT(1416)  = ~\3851GAT(1392)  & ~\3850GAT(1379) ,
  \2007GAT(604)  = ~\1831GAT(540)  & ~\1951GAT(576) ,
  \1829GAT(538)  = ~\1767GAT(499)  & ~\1720GAT(482) ,
  \1763GAT(500)  = ~\549GAT(285)  & ~\1717GAT(483) ,
  \[20]  = ~\6186GAT(2396)  & ~\6185GAT(2395) ,
  \5460GAT(2078)  = ~\1065GAT(113)  & ~\5404GAT(2052) ,
  \[21]  = ~\6196GAT(2401)  & ~\6195GAT(2400) ,
  \2342GAT(726)  = ~\2301GAT(708)  & ~\2248GAT(691) ,
  \3632GAT(1288)  = ~\3516GAT(1237)  & ~\3574GAT(1265) ,
  \6068GAT(2343)  = ~\6040GAT(2335)  & ~\6011GAT(2319) ,
  \[22]  = ~\6206GAT(2406)  & ~\6205GAT(2405) ,
  \1167GAT(79)  = \273GAT(16)  & \222GAT(13) ,
  \1152GAT(84)  = \460GAT(27)  & \205GAT(12) ,
  \1821GAT(484)  = ~\1759GAT(470)  & ~\1624GAT(408) ,
  \[23]  = ~\6216GAT(2411)  & ~\6215GAT(2410) ,
  \2043GAT(620)  = ~\2009GAT(602)  & ~\2008GAT(599) ,
  \3667GAT(1320)  = ~\3491GAT(1249)  & ~\3612GAT(1293) ,
  \3874GAT(1372)  = ~\3805GAT(1350)  & ~\3804GAT(1349) ,
  \1335GAT(296)  = ~\879GAT(175) ,
  \1876GAT(513)  = ~\1803GAT(490)  & ~\1668GAT(429) ,
  \1397GAT(306)  = ~\1363GAT(289)  & ~\1215GAT(63) ,
  \[24]  = ~\6226GAT(2416)  & ~\6225GAT(2415) ,
  \[25]  = ~\6236GAT(2421)  & ~\6235GAT(2420) ,
  \[26]  = ~\6246GAT(2426)  & ~\6245GAT(2425) ,
  \1702GAT(451)  = ~\1660GAT(431)  & ~\1606GAT(414) ,
  \[27]  = ~\6256GAT(2431)  & ~\6255GAT(2430) ,
  \5989GAT(2310)  = ~\828GAT(192)  & ~\5950GAT(2292) ,
  \2902GAT(973)  = ~\2852GAT(941)  & ~\2851GAT(933) ,
  \2668GAT(876)  = ~\2513GAT(803)  & ~\2623GAT(851) ,
  \5434GAT(2081)  = ~\774GAT(210)  & ~\5380GAT(2049) ,
  \[28]  = ~\6266GAT(2436)  & ~\6265GAT(2435) ,
  \2305GAT(707)  = ~\2196GAT(656)  & ~\2251GAT(690) ,
  \1820GAT(486)  = ~\1221GAT(61)  & ~\1759GAT(470) ,
  \[29]  = ~\6276GAT(2441)  & ~\6275GAT(2440) ,
  \2789GAT(913)  = ~\2727GAT(899)  & ~\2675GAT(863) ,
  \2006GAT(601)  = ~\1951GAT(576)  & ~\1905GAT(559) ,
  \1158GAT(82)  = \494GAT(29)  & \205GAT(12) ,
  \2181GAT(665)  = ~\2109GAT(634)  & ~\1971GAT(571) ,
  \4395GAT(1597)  = ~\4344GAT(1585)  & ~\4167GAT(1496) ,
  \2341GAT(733)  = ~\2186GAT(662)  & ~\2297GAT(709) ,
  \5399GAT(2043)  = ~\5339GAT(2019)  & ~\5280GAT(1986) ,
  \4377GAT(1603)  = ~\4328GAT(1586)  & ~\4327GAT(1581) ,
  \2488GAT(818)  = ~\2422GAT(780)  & ~\2277GAT(714) ,
  \1155GAT(83)  = \477GAT(28)  & \205GAT(12) ,
  \1704GAT(449)  = ~\1664GAT(430)  & ~\1609GAT(413) ,
  \5594GAT(2113)  = ~\5531GAT(2104)  & ~\5473GAT(2059) ,
  \6217GAT(2409)  = ~\6211GAT(2407)  & ~\5962GAT(2280) ,
  \3718GAT(1337)  = ~\3671GAT(1318)  & ~\3670GAT(1308) ,
  \[30]  = ~\6281GAT(2442)  & ~\5602GAT(2110) ,
  \948GAT(152)  = \392GAT(23)  & \137GAT(8) ,
  \3166GAT(1098)  = ~\801GAT(201)  & ~\3099GAT(1064) ,
  \2966GAT(989)  = ~\2908GAT(970)  & ~\2861GAT(930) ,
  \[31]  = ~\6286GAT(2446)  & ~\6285GAT(2445) ,
  \3305GAT(1138)  = ~\1092GAT(104)  & ~\3245GAT(1113) ,
  \4365GAT(1606)  = ~\4319GAT(1588)  & ~\4318GAT(1583) ,
  \2180GAT(667)  = ~\840GAT(188)  & ~\2109GAT(634) ,
  \4716GAT(1762)  = ~\4662GAT(1743)  & ~\4604GAT(1715) ,
  \4825GAT(1819)  = ~\672GAT(244)  & ~\4766GAT(1792) ,
  \1396GAT(307)  = ~\1359GAT(290) ,
  \3592GAT(1259)  = ~\3536GAT(1230)  & ~\3356GAT(1152) ,
  \4572GAT(1674)  = ~\4503GAT(1661)  & ~\4335GAT(1578) ,
  \5560GAT(2124)  = ~\5495GAT(2099)  & ~\5498GAT(2098) ,
  \840GAT(188)  = \324GAT(19)  & \103GAT(6) ,
  \3199GAT(1072)  = ~\3132GAT(1053)  & ~\3131GAT(1052) ,
  \972GAT(144)  = \528GAT(31)  & \137GAT(8) ,
  \2395GAT(750)  = ~\2349GAT(725)  & ~\2348GAT(720) ,
  \2828GAT(954)  = ~\2761GAT(921)  & ~\2611GAT(854) ,
  \1738GAT(476)  = ~\1701GAT(454)  & ~\1700GAT(453) ,
  \5575GAT(2119)  = ~\5510GAT(2107)  & ~\5339GAT(2019) ,
  \5069GAT(1919)  = ~\5013GAT(1900)  & ~\4953GAT(1871) ,
  \1926GAT(552)  = ~\1870GAT(518)  & ~\1869GAT(514) ,
  \3079GAT(1069)  = ~\561GAT(281)  & ~\3028GAT(1050) ,
  \6089GAT(2353)  = ~\6064GAT(2346)  & ~\6037GAT(2332) ,
  \3734GAT(1331)  = ~\3681GAT(1312)  & ~\3638GAT(1283) ,
  \5607GAT(2166)  = ~\582GAT(274)  & ~\5540GAT(2135) ,
  \6031GAT(2314)  = ~\5956GAT(2282)  & ~\5996GAT(2300) ,
  \1703GAT(452)  = ~\1548GAT(381)  & ~\1660GAT(431) ,
  \2005GAT(605)  = ~\1826GAT(543)  & ~\1947GAT(577) ,
  \5193GAT(1973)  = ~\771GAT(211)  & ~\5130GAT(1952) ,
  \4394GAT(1609)  = ~\1200GAT(68)  & ~\4344GAT(1585) ,
  \816GAT(196)  = \460GAT(27)  & \86GAT(5) ,
  \4432GAT(1633)  = ~\4373GAT(1615)  & ~\4372GAT(1605) ,
  \4668GAT(1736)  = ~\4612GAT(1713)  & ~\4611GAT(1712) ,
  \4034GAT(1449)  = ~\3986GAT(1429)  & ~\3989GAT(1428) ,
  \1660GAT(431)  = ~\1548GAT(381)  & ~\1606GAT(414) ,
  \2223GAT(700)  = \[3] ,
  \5085GAT(1914)  = ~\5031GAT(1896)  & ~\5030GAT(1891) ,
  \1395GAT(308)  = ~\1359GAT(290)  & ~\1167GAT(79) ,
  \3675GAT(1316)  = ~\3511GAT(1240)  & ~\3628GAT(1289) ,
  \4754GAT(1750)  = ~\4698GAT(1727)  & ~\4701GAT(1726) ,
  \1197GAT(69)  = \443GAT(26)  & \222GAT(13) ,
  \1005GAT(133)  = \443GAT(26)  & \154GAT(9) ,
  \3804GAT(1349)  = ~\3742GAT(1328)  & ~\3690GAT(1300) ,
  \4420GAT(1636)  = ~\4364GAT(1617)  & ~\4363GAT(1607) ,
  \672GAT(244)  = \460GAT(27)  & \35GAT(2) ,
  \4450GAT(1627)  = ~\4389GAT(1611)  & ~\4232GAT(1520) ,
  \4921GAT(1843)  = ~\1011GAT(131)  & ~\4854GAT(1815) ,
  \3603GAT(1256)  = ~\3476GAT(1196)  & ~\3548GAT(1217) ,
  \4216GAT(1526)  = ~\4079GAT(1481)  & ~\4146GAT(1503) ,
  \3955GAT(1441)  = ~\3837GAT(1397)  & ~\3902GAT(1419) ,
  \1880GAT(512)  = ~\1077GAT(109)  & ~\1807GAT(489) ,
  \558GAT(282)  = \358GAT(21)  & \1GAT(0) ,
  \5552GAT(2127)  = ~\5489GAT(2109)  & ~\5431GAT(2073) ,
  \5446GAT(2069)  = ~\5389GAT(2047)  & ~\5392GAT(2046) ,
  \5797GAT(2234)  = ~\777GAT(209)  & ~\5743GAT(2211) ,
  \4866GAT(1802)  = ~\4802GAT(1781)  & ~\4805GAT(1780) ,
  \2359GAT(717)  = ~\2322GAT(703)  & ~\2145GAT(623) ,
  \2587GAT(826)  = ~\2464GAT(768)  & ~\2539GAT(786) ,
  \6237GAT(2419)  = ~\6231GAT(2417)  & ~\5873GAT(2241) ,
  \2260GAT(687)  = ~\2211GAT(647)  & ~\2214GAT(644) ,
  \1462GAT(358)  = ~\738GAT(222)  & ~\1413GAT(343) ,
  \3809GAT(1356)  = ~\1146GAT(86)  & ~\3748GAT(1325) ,
  \3608GAT(1294)  = ~\3486GAT(1251)  & ~\3556GAT(1273) ,
  \1101GAT(101)  = \443GAT(26)  & \188GAT(11) ,
  \5354GAT(2014)  = ~\5292GAT(1998)  & ~\5109GAT(1906) ,
  \5267GAT(1991)  = ~\5136GAT(1942)  & ~\5200GAT(1965) ,
  \1826GAT(543)  = ~\1763GAT(500)  & ~\1628GAT(439) ,
  \5764GAT(2209)  = ~\1020GAT(128)  & ~\5706GAT(2174) ,
  \3506GAT(1243)  = ~\3437GAT(1211)  & ~\3284GAT(1143) ,
  \4900GAT(1846)  = ~\768GAT(212)  & ~\4833GAT(1817) ,
  \621GAT(261)  = \443GAT(26)  & \18GAT(1) ,
  \1543GAT(384)  = ~\1474GAT(355)  & ~\1339GAT(295) ,
  \1478GAT(354)  = ~\930GAT(158)  & ~\1425GAT(339) ,
  \3212GAT(1127)  = ~\3146GAT(1106)  & ~\3145GAT(1094) ,
  \2426GAT(779)  = ~\699GAT(235)  & ~\2371GAT(760) ,
  \2358GAT(721)  = ~\1227GAT(59)  & ~\2322GAT(703) ,
  \873GAT(177)  = \511GAT(30)  & \103GAT(6) ,
  \1881GAT(510)  = ~\1807GAT(489)  & ~\1672GAT(428) ,
  \753GAT(217)  = \375GAT(22)  & \69GAT(4) ,
  \1753GAT(471)  = ~\1711GAT(444)  & ~\1710GAT(443) ,
  \4913GAT(1831)  = ~\4850GAT(1808)  & ~\4849GAT(1807) ,
  \2004GAT(603)  = ~\1947GAT(577)  & ~\1902GAT(560) ,
  \6046GAT(2330)  = ~\6014GAT(2322)  & ~\5898GAT(2268) ,
  \4598GAT(1719)  = ~\4540GAT(1695)  & ~\4539GAT(1684) ,
  \1394GAT(309)  = ~\1355GAT(291) ,
  \6240GAT(2423)  = \[25] ,
  \6250GAT(2428)  = \[26] ,
  \1588GAT(420)  = ~\1522GAT(398)  & ~\1521GAT(397) ,
  \1401GAT(347)  = ~\1372GAT(331)  & ~\1371GAT(332) ,
  \3124GAT(1055)  = ~\3063GAT(1043)  & ~\3062GAT(1038) ,
  \2753GAT(923)  = ~\654GAT(250)  & ~\2700GAT(904) ,
  \4358GAT(1620)  = ~\4185GAT(1546)  & ~\4302GAT(1592) ,
  \5021GAT(1893)  = ~\4959GAT(1869)  & ~\4904GAT(1835) ,
  \1542GAT(386)  = ~\882GAT(174)  & ~\1474GAT(355) ,
  \2864GAT(929)  = ~\2791GAT(912)  & ~\2794GAT(911) ,
  \5919GAT(2261)  = ~\5867GAT(2243)  & ~\5870GAT(2242) ,
  \2277GAT(714)  = ~\2161GAT(677)  & ~\2230GAT(697) ,
  \5685GAT(2181)  = ~\5629GAT(2151)  & ~\5628GAT(2150) ,
  \5808GAT(2223)  = ~\5755GAT(2202)  & ~\5697GAT(2178) ,
  \2513GAT(803)  = ~\2442GAT(775)  & ~\2297GAT(709) ,
  \1017GAT(129)  = \511GAT(30)  & \154GAT(9) ,
  \6061GAT(2344)  = ~\6036GAT(2336)  & ~\6035GAT(2333) ,
  \5895GAT(2269)  = ~\5845GAT(2256)  & ~\5844GAT(2251) ,
  \4012GAT(1468)  = ~\3842GAT(1395)  & ~\3959GAT(1440) ,
  \4161GAT(1498)  = ~\4094GAT(1487)  & ~\3938GAT(1406) ,
  \591GAT(271)  = \273GAT(16)  & \18GAT(1) ,
  \5250GAT(2005)  = ~\675GAT(243)  & ~\5184GAT(1975) ,
  \1083GAT(107)  = \341GAT(20)  & \188GAT(11) ,
  \3637GAT(1287)  = ~\3521GAT(1234)  & ~\3577GAT(1264) ,
  \2257GAT(688)  = ~\2210GAT(649)  & ~\2209GAT(645) ,
  \1815GAT(487)  = ~\1173GAT(77)  & ~\1756GAT(469) ,
  \6056GAT(2326)  = ~\6026GAT(2315)  & ~\5993GAT(2301) ,
  \1191GAT(71)  = \409GAT(24)  & \222GAT(13) ,
  \5727GAT(2167)  = ~\5671GAT(2137)  & ~\5670GAT(2136) ,
  \5035GAT(1889)  = ~\4973GAT(1877)  & ~\4972GAT(1865) ,
  \702GAT(234)  = \358GAT(21)  & \52GAT(3) ,
  \4529GAT(1686)  = ~\4466GAT(1667)  & ~\4408GAT(1642) ,
  \1825GAT(544)  = ~\549GAT(285)  & ~\1763GAT(500) ,
  \810GAT(198)  = \426GAT(25)  & \86GAT(5) ,
  \1194GAT(70)  = \426GAT(25)  & \222GAT(13) ,
  \5480GAT(2105)  = ~\5426GAT(2084)  & ~\5425GAT(2077) ,
  \4748GAT(1752)  = ~\4692GAT(1739)  & ~\4515GAT(1649) ,
  \870GAT(178)  = \494GAT(29)  & \103GAT(6) ,
  \1014GAT(130)  = \494GAT(29)  & \154GAT(9) ,
  \2502GAT(811)  = ~\795GAT(203)  & ~\2434GAT(777) ,
  \5047GAT(1895)  = ~\1110GAT(98)  & ~\4986GAT(1859) ,
  \5353GAT(2030)  = ~\1161GAT(81)  & ~\5292GAT(1998) ,
  \2718GAT(896)  = ~\2670GAT(874)  & ~\2669GAT(867) ,
  \3676GAT(1304)  = ~\3632GAT(1288)  & ~\3574GAT(1265) ,
  \5608GAT(2165)  = ~\5540GAT(2135)  & ~\5366GAT(2058) ,
  \2586GAT(825)  = ~\2539GAT(786)  & ~\2467GAT(767) ,
  \3248GAT(1121)  = ~\1140GAT(88)  & ~\3199GAT(1072) ,
  \3668GAT(1309)  = ~\3616GAT(1292)  & ~\3562GAT(1271) ,
  \2512GAT(805)  = ~\891GAT(171)  & ~\2442GAT(775) ,
  \1331GAT(297)  = ~\831GAT(191) ,
  \795GAT(203)  = \341GAT(20)  & \86GAT(5) ,
  \4787GAT(1786)  = ~\4727GAT(1759)  & ~\4730GAT(1758) ,
  \2101GAT(636)  = ~\744GAT(220)  & ~\2049GAT(618) ,
  \2236GAT(695)  = ~\2175GAT(670)  & ~\2174GAT(663) ,
  \6151GAT(2377)  = ~\6147GAT(2374)  & ~\6135GAT(2369) ,
  \1929GAT(551)  = ~\1875GAT(515)  & ~\1874GAT(511) ,
  \3515GAT(1239)  = ~\900GAT(168)  & ~\3445GAT(1209) ,
  \6267GAT(2434)  = ~\6261GAT(2432)  & ~\5721GAT(2170) ,
  \5344GAT(2018)  = ~\5215GAT(1960)  & ~\5283GAT(1985) ,
  \3841GAT(1396)  = ~\711GAT(231)  & ~\3772GAT(1362) ,
  \1750GAT(472)  = ~\1709GAT(446)  & ~\1708GAT(445) ,
  \1824GAT(541)  = ~\1763GAT(500)  & ~\1717GAT(483) ,
  \6141GAT(2373)  = ~\6138GAT(2372) ,
  \5734GAT(2213)  = ~\5613GAT(2163)  & ~\5676GAT(2185) ,
  \5709GAT(2189)  = ~\1068GAT(112)  & ~\5651GAT(2142) ,
  \2785GAT(915)  = ~\1038GAT(122)  & ~\2724GAT(894) ,
  \1618GAT(410)  = ~\1572GAT(368)  & ~\1571GAT(367) ,
  \2913GAT(969)  = ~\2791GAT(912)  & ~\2864GAT(929) ,
  \2309GAT(706)  = ~\2201GAT(653)  & ~\2254GAT(689) ,
  \5861GAT(2255)  = ~\924GAT(160)  & ~\5810GAT(2222) ,
  \2398GAT(754)  = ~\1131GAT(91)  & ~\2350GAT(719) ,
  \4526GAT(1700)  = ~\4462GAT(1668)  & ~\4294GAT(1594) ,
  \1541GAT(385)  = ~\1474GAT(355)  & ~\1422GAT(340) ,
  \4049GAT(1444)  = ~\4001GAT(1433)  & ~\3821GAT(1344) ,
  \3091GAT(1066)  = ~\705GAT(233)  & ~\3037GAT(1047) ,
  \4677GAT(1734)  = ~\4616GAT(1724)  & ~\4435GAT(1632) ,
  \4298GAT(1593)  = ~\4180GAT(1548)  & ~\4245GAT(1568) ,
  \4122GAT(1513)  = ~\714GAT(230)  & ~\4061GAT(1488) ,
  \6018GAT(2318)  = ~\5984GAT(2311)  & ~\5947GAT(2284) ,
  \4508GAT(1660)  = ~\1104GAT(100)  & ~\4444GAT(1641) ,
  \5240GAT(2009)  = ~\579GAT(275)  & ~\5176GAT(1977) ,
  \4318GAT(1583)  = ~\4260GAT(1562)  & ~\4208GAT(1528) ,
  \4110GAT(1516)  = ~\570GAT(278)  & ~\4052GAT(1491) ,
  \6255GAT(2430)  = ~\6251GAT(2427)  & ~\5879GAT(2238) ,
  \5426GAT(2084)  = ~\5241GAT(2008)  & ~\5366GAT(2058) ,
  \3190GAT(1076)  = ~\3120GAT(1059)  & ~\3119GAT(1057) ,
  \5471GAT(2060)  = ~\5416GAT(2038)  & ~\5357GAT(2013) ,
  \3527GAT(1224)  = ~\3455GAT(1203)  & ~\3458GAT(1202) ,
  \6190GAT(2398)  = \[20] ,
  \5829GAT(2216)  = ~\5776GAT(2195)  & ~\5718GAT(2171) ,
  \3917GAT(1413)  = ~\3862GAT(1386)  & ~\3865GAT(1376) ,
  \1116GAT(96)  = \528GAT(31)  & \188GAT(11) ,
  \2281GAT(713)  = ~\2166GAT(674)  & ~\2233GAT(696) ,
  \2503GAT(809)  = ~\2434GAT(777)  & ~\2289GAT(711) ,
  \2061GAT(614)  = ~\2021GAT(590)  & ~\2020GAT(587) ,
  \3037GAT(1047)  = ~\2994GAT(1028)  & ~\2993GAT(1020) ,
  \2117GAT(632)  = ~\936GAT(156)  & ~\2061GAT(614) ,
  \3185GAT(1077)  = ~\3115GAT(1060)  & ~\3055GAT(1039) ,
  \3075GAT(1034)  = ~\2977GAT(986)  & ~\3022GAT(1005) ,
  \5930GAT(2295)  = ~\5882GAT(2276)  & ~\5730GAT(2214) ,
  \6101GAT(2348)  = ~\6076GAT(2340)  & ~\6049GAT(2329) ,
  \2527GAT(796)  = ~\1035GAT(123)  & ~\2454GAT(772) ,
  \3067GAT(1036)  = ~\3015GAT(1013)  & ~\3014GAT(1008) ,
  \2230GAT(697)  = ~\2165GAT(676)  & ~\2164GAT(669) ,
  \2912GAT(968)  = ~\2864GAT(929)  & ~\2794GAT(911) ,
  \2497GAT(814)  = ~\747GAT(219)  & ~\2430GAT(778) ,
  \2349GAT(725)  = ~\2206GAT(650)  & ~\2313GAT(705) ,
  \1571GAT(367)  = ~\1498GAT(349)  & ~\1440GAT(334) ,
  \4211GAT(1527)  = ~\4140GAT(1505)  & ~\4143GAT(1504) ,
  \906GAT(166)  = \426GAT(25)  & \120GAT(7) ,
  \1119GAT(95)  = \273GAT(16)  & \205GAT(12) ,
  \2573GAT(831)  = ~\2522GAT(799)  & ~\2521GAT(790) ,
  \2174GAT(663)  = ~\2105GAT(635)  & ~\2052GAT(617) ,
  \5759GAT(2200)  = ~\5700GAT(2177)  & ~\5642GAT(2146) ,
  \3000GAT(1023)  = ~\2838GAT(948)  & ~\2950GAT(996) ,
  \4863GAT(1803)  = ~\4801GAT(1794)  & ~\4800GAT(1782) ,
  \3620GAT(1291)  = ~\3501GAT(1245)  & ~\3565GAT(1269) ,
  \2470GAT(766)  = ~\2404GAT(748)  & ~\2407GAT(747) ,
  \5331GAT(2022)  = ~\5271GAT(2001)  & ~\5206GAT(1962) ,
  \1518GAT(399)  = ~\1454GAT(360)  & ~\1319GAT(300) ,
  \4621GAT(1723)  = ~\1008GAT(132)  & ~\4566GAT(1689) ,
  \4812GAT(1777)  = ~\4754GAT(1750)  & ~\4701GAT(1726) ,
  \1113GAT(97)  = \511GAT(30)  & \188GAT(11) ,
  \1110GAT(98)  = \494GAT(29)  & \188GAT(11) ,
  \1585GAT(421)  = ~\1517GAT(401)  & ~\1516GAT(400) ,
  \2009GAT(602)  = ~\1836GAT(537)  & ~\1955GAT(575) ,
  \4859GAT(1814)  = ~\1059GAT(115)  & ~\4796GAT(1796) ,
  \2749GAT(924)  = ~\606GAT(266)  & ~\2697GAT(905) ,
  \3872GAT(1373)  = ~\3800GAT(1351)  & ~\3739GAT(1329) ,
  \5221GAT(1958)  = ~\5157GAT(1935)  & ~\5160GAT(1934) ,
  \4405GAT(1643)  = ~\4354GAT(1622)  & ~\4353GAT(1614) ,
  \1122GAT(94)  = \290GAT(17)  & \205GAT(12) ,
  \5878GAT(2240)  = ~\5770GAT(2197)  & ~\5825GAT(2218) ,
  \3227GAT(1122)  = ~\3171GAT(1095)  & ~\3170GAT(1082) ,
  \2794GAT(911)  = ~\2732GAT(897)  & ~\2731GAT(893) ,
  \4950GAT(1873)  = ~\4890GAT(1850)  & ~\4889GAT(1840) ,
  \3325GAT(1168)  = ~\3268GAT(1147)  & ~\3215GAT(1126) ,
  \6166GAT(2386)  = ~\6157GAT(2379)  & ~\6161GAT(2382) ,
  \5990GAT(2302)  = ~\5950GAT(2292)  & ~\5804GAT(2225) ,
  \1020GAT(128)  = \528GAT(31)  & \154GAT(9) ,
  \1080GAT(108)  = \324GAT(19)  & \188GAT(11) ,
  \2254GAT(689)  = ~\2205GAT(652)  & ~\2204GAT(646) ,
  \3215GAT(1126)  = ~\3151GAT(1104)  & ~\3150GAT(1091) ,
  \915GAT(163)  = \477GAT(28)  & \120GAT(7) ,
  \2348GAT(720)  = ~\2313GAT(705)  & ~\2257GAT(688) ,
  \3541GAT(1228)  = ~\1191GAT(71)  & ~\3470GAT(1206) ,
  \3476GAT(1196)  = ~\3413GAT(1185)  & ~\3260GAT(1109) ,
  \5749GAT(2204)  = ~\5688GAT(2191)  & ~\5501GAT(2097) ,
  \3131GAT(1052)  = ~\3070GAT(1035)  & ~\3019GAT(1006) ,
  \5464GAT(2063)  = ~\5409GAT(2051)  & ~\5408GAT(2041) ,
  \4487GAT(1662)  = ~\861GAT(181)  & ~\4423GAT(1645) ,
  \5194GAT(1967)  = ~\5130GAT(1952)  & ~\4959GAT(1869) ,
  \5136GAT(1942)  = ~\5076GAT(1925)  & ~\4907GAT(1834) ,
  \1128GAT(92)  = \324GAT(19)  & \205GAT(12) ,
  \5065GAT(1921)  = ~\5005GAT(1902)  & ~\4947GAT(1875) ,
  \3257GAT(1110)  = ~\3207GAT(1078)  & ~\3206GAT(1071) ,
  \2049GAT(618)  = ~\2013GAT(598)  & ~\2012GAT(595) ,
  \5280GAT(1986)  = ~\5214GAT(1971)  & ~\5213GAT(1961) ,
  \6245GAT(2425)  = ~\6241GAT(2422)  & ~\5925GAT(2258) ,
  \1787GAT(494)  = ~\837GAT(189)  & ~\1735GAT(477) ,
  \5531GAT(2104)  = ~\1212GAT(64)  & ~\5473GAT(2059) ,
  \4696GAT(1728)  = ~\4637GAT(1718)  & ~\4584GAT(1669) ,
  \5124GAT(1946)  = ~\5070GAT(1927)  & ~\5069GAT(1919) ,
  \4613GAT(1711)  = ~\4562GAT(1678)  & ~\4561GAT(1677) ,
  \4998GAT(1856)  = ~\4942GAT(1837)  & ~\4941GAT(1823) ,
  \813GAT(197)  = \443GAT(26)  & \86GAT(5) ,
  \1399GAT(304)  = ~\1367GAT(288)  & ~\1263GAT(47) ,
  \5587GAT(2114)  = ~\5527GAT(2089)  & ~\5526GAT(2088) ,
  \4871GAT(1801)  = ~\4748GAT(1752)  & ~\4808GAT(1779) ,
  \4544GAT(1683)  = ~\4478GAT(1664)  & ~\4417GAT(1637) ,
  \1125GAT(93)  = \307GAT(18)  & \205GAT(12) ,
  \5971GAT(2309)  = \[14] ,
  \2176GAT(668)  = ~\2105GAT(635)  & ~\1967GAT(572) ,
  \3556GAT(1273)  = ~\3490GAT(1250)  & ~\3489GAT(1235) ,
  \2877GAT(983)  = \[5] ,
  \4709GAT(1775)  = ~\4526GAT(1700)  & ~\4646GAT(1747) ,
  \2968GAT(988)  = ~\2913GAT(969)  & ~\2912GAT(968) ,
  \2008GAT(599)  = ~\1955GAT(575)  & ~\1908GAT(558) ,
  \5343GAT(2017)  = ~\5283GAT(1985)  & ~\5218GAT(1959) ,
  \4017GAT(1454)  = ~\3971GAT(1437)  & ~\3914GAT(1414) ,
  \5670GAT(2136)  = ~\5602GAT(2110)  & ~\1308GAT(32) ,
  \615GAT(263)  = \409GAT(24)  & \18GAT(1) ,
  \6023GAT(2316)  = ~\5989GAT(2310)  & ~\5988GAT(2303) ,
  \2570GAT(832)  = ~\2517GAT(802)  & ~\2516GAT(792) ,
  \5886GAT(2275)  = ~\633GAT(257)  & ~\5837GAT(2252) ,
  \2517GAT(802)  = ~\939GAT(155)  & ~\2446GAT(774) ,
  \909GAT(165)  = \443GAT(26)  & \120GAT(7) ,
  \2486GAT(810)  = ~\2422GAT(780)  & ~\2368GAT(761) ,
  \2870GAT(926)  = ~\2802GAT(909)  & ~\2801GAT(908) ,
  \1023GAT(127)  = \273GAT(16)  & \171GAT(10) ,
  \6064GAT(2346)  = ~\636GAT(256)  & ~\6037GAT(2332) ,
  \1831GAT(540)  = ~\1767GAT(499)  & ~\1632GAT(438) ,
  \3836GAT(1398)  = ~\663GAT(247)  & ~\3768GAT(1363) ,
  \1732GAT(478)  = ~\1697GAT(458)  & ~\1696GAT(457) ,
  \5693GAT(2190)  = ~\873GAT(177)  & ~\5633GAT(2160) ,
  \2175GAT(670)  = ~\792GAT(204)  & ~\2105GAT(635) ,
  \1131GAT(91)  = \341GAT(20)  & \205GAT(12) ,
  \5867GAT(2243)  = ~\5813GAT(2233)  & ~\5645GAT(2145) ,
  \5081GAT(1924)  = ~\867GAT(179)  & ~\5026GAT(1897) ,
  \1640GAT(436)  = ~\1523GAT(396)  & ~\1591GAT(419) ,
  \5438GAT(2072)  = ~\5383GAT(2054)  & ~\5324GAT(2023) ,
  \1104GAT(100)  = \460GAT(27)  & \188GAT(11) ,
  \1573GAT(366)  = ~\1498GAT(349)  & ~\1363GAT(289) ,
  \4829GAT(1818)  = ~\720GAT(228)  & ~\4769GAT(1791) ,
  \1134GAT(90)  = \358GAT(21)  & \205GAT(12) ,
  \5324GAT(2023)  = ~\5267GAT(1991)  & ~\5266GAT(1990) ,
  \6070GAT(2342)  = ~\6040GAT(2335)  & ~\5941GAT(2287) ,
  \1398GAT(305)  = ~\1363GAT(289) ,
  \2487GAT(819)  = ~\651GAT(251)  & ~\2422GAT(780) ,
  \3337GAT(1158)  = ~\3292GAT(1141)  & ~\3233GAT(1118) ,
  \5612GAT(2164)  = ~\630GAT(258)  & ~\5544GAT(2134) ,
  \2501GAT(801)  = ~\2434GAT(777)  & ~\2377GAT(758) ,
  \6186GAT(2396)  = ~\6177GAT(2389)  & ~\6181GAT(2392) ,
  \6011GAT(2319)  = ~\5980GAT(2306)  & ~\5979GAT(2305) ,
  \3681GAT(1312)  = ~\999GAT(135)  & ~\3638GAT(1283) ,
  \4928GAT(1827)  = ~\4860GAT(1804)  & ~\4863GAT(1803) ,
  \2521GAT(790)  = ~\2450GAT(773)  & ~\2389GAT(753) ,
  \6128GAT(2365)  = ~\6114GAT(2359)  & ~\6094GAT(2351) ,
  \5348GAT(2032)  = ~\1113GAT(97)  & ~\5289GAT(1982) ,
  \4099GAT(1485)  = ~\1197GAT(69)  & ~\4043GAT(1457) ,
  \2967GAT(992)  = ~\2858GAT(936)  & ~\2908GAT(970) ,
  \3673GAT(1317)  = ~\3506GAT(1243)  & ~\3624GAT(1290) ,
  \3851GAT(1392)  = ~\807GAT(199)  & ~\3780GAT(1360) ,
  \4885GAT(1852)  = ~\624GAT(260)  & ~\4821GAT(1820) ,
  \5947GAT(2284)  = ~\5903GAT(2267)  & ~\5902GAT(2266) ,
  \4895GAT(1848)  = ~\720GAT(228)  & ~\4829GAT(1818) ,
  \1092GAT(104)  = \392GAT(23)  & \188GAT(11) ,
  \1819GAT(485)  = ~\1759GAT(470)  & ~\1714GAT(440) ,
  \2873GAT(932)  = ~\1233GAT(57)  & ~\2803GAT(907) ,
  \2663GAT(873)  = ~\2615GAT(853)  & ~\2564GAT(834) ,
  \5721GAT(2170)  = ~\5660GAT(2140)  & ~\5663GAT(2139) ,
  \2995GAT(1018)  = ~\2942GAT(998)  & ~\2890GAT(978) ,
  \552GAT(284)  = \324GAT(19)  & \1GAT(0) ,
  \2662GAT(882)  = ~\2498GAT(812)  & ~\2611GAT(854) ,
  \3815GAT(1346)  = ~\3751GAT(1335)  & ~\3598GAT(1257) ,
  \4530GAT(1699)  = ~\621GAT(261)  & ~\4466GAT(1667) ,
  \5713GAT(2173)  = ~\5654GAT(2158)  & ~\5587GAT(2114) ,
  \6085GAT(2355)  = ~\588GAT(272)  & ~\6061GAT(2344) ,
  \2522GAT(799)  = ~\987GAT(139)  & ~\2450GAT(773) ,
  \4040GAT(1446)  = ~\3997GAT(1426)  & ~\3996GAT(1425) ,
  \5188GAT(1974)  = ~\723GAT(227)  & ~\5127GAT(1944) ,
  \2357GAT(718)  = ~\2322GAT(703)  & ~\2266GAT(684) ,
  \5218GAT(1959)  = ~\5156GAT(1949)  & ~\5155GAT(1936) ,
  \1668GAT(429)  = ~\1558GAT(375)  & ~\1612GAT(412) ,
  \1086GAT(106)  = \358GAT(21)  & \188GAT(11) ,
  \2179GAT(660)  = ~\2109GAT(634)  & ~\2055GAT(616) ,
  \4946GAT(1876)  = \[11] ,
  \5304GAT(1978)  = ~\5236GAT(1953)  & ~\1305GAT(33) ,
  \1572GAT(368)  = ~\1170GAT(78)  & ~\1498GAT(349) ,
  \2076GAT(611)  = ~\1176GAT(76)  & ~\2030GAT(578) ,
  \2639GAT(844)  = ~\2582GAT(827)  & ~\2536GAT(787) ,
  \2233GAT(696)  = ~\2170GAT(673)  & ~\2169GAT(666) ,
  \3509GAT(1229)  = ~\3441GAT(1210)  & ~\3383GAT(1187) ,
  \4143GAT(1504)  = ~\4078GAT(1492)  & ~\4077GAT(1482) ,
  \2703GAT(903)  = ~\2660GAT(884)  & ~\2659GAT(877) ,
  \6197GAT(2399)  = ~\6191GAT(2397)  & ~\6026GAT(2315) ,
  \3805GAT(1350)  = ~\3687GAT(1301)  & ~\3742GAT(1328) ,
  \4680GAT(1733)  = ~\4621GAT(1723)  & ~\4620GAT(1710) ,
  \4389GAT(1611)  = ~\1152GAT(84)  & ~\4341GAT(1575) ,
  \4984GAT(1860)  = ~\4928GAT(1827)  & ~\4863GAT(1803) ,
  \4043GAT(1457)  = ~\1197GAT(69)  & ~\3998GAT(1424) ,
  \1830GAT(542)  = ~\597GAT(269)  & ~\1767GAT(499) ,
  \2715GAT(898)  = ~\2668GAT(876)  & ~\2667GAT(869) ,
  \1050GAT(118)  = \426GAT(25)  & \171GAT(10) ,
  \1400GAT(303)  = ~\1367GAT(288) ,
  \5494GAT(2108)  = ~\774GAT(210)  & ~\5434GAT(2081) ,
  \2222GAT(642)  = ~\2082GAT(606)  & ~\2145GAT(623) ,
  \2345GAT(729)  = ~\2196GAT(656)  & ~\2305GAT(707) ,
  \5234GAT(1954)  = ~\5172GAT(1945)  & ~\5115GAT(1903) ,
  \6082GAT(2337)  = ~\6057GAT(2327)  & ~\6056GAT(2326) ,
  \4175GAT(1550)  = ~\4110GAT(1516)  & ~\3947GAT(1443) ,
  \5289GAT(1982)  = ~\5226GAT(1957)  & ~\5225GAT(1956) ,
  \5935GAT(2293)  = ~\5886GAT(2275)  & ~\5734GAT(2213) ,
  \1694GAT(459)  = ~\1644GAT(435)  & ~\1594GAT(418) ,
  \2536GAT(787)  = ~\2463GAT(770)  & ~\2462GAT(769) ,
  \4264GAT(1560)  = ~\4211GAT(1527)  & ~\4143GAT(1504) ,
  \5873GAT(2241)  = ~\5819GAT(2220)  & ~\5822GAT(2219) ,
  \3604GAT(1295)  = ~\3481GAT(1253)  & ~\3553GAT(1274) ,
  \3165GAT(1083)  = ~\3099GAT(1064)  & ~\3043GAT(1044) ,
  \3582GAT(1263)  = ~\3455GAT(1203)  & ~\3527GAT(1224) ,
  \6196GAT(2401)  = ~\6187GAT(2394)  & ~\6191GAT(2397) ,
  \5101GAT(1909)  = ~\5047GAT(1895)  & ~\4986GAT(1859) ,
  \798GAT(202)  = \358GAT(21)  & \86GAT(5) ,
  \3147GAT(1105)  = ~\3083GAT(1068)  & ~\2930GAT(1001) ,
  \1146GAT(86)  = \426GAT(25)  & \205GAT(12) ,
  \2797GAT(910)  = ~\2733GAT(892)  & ~\2736GAT(891) ,
  \3986GAT(1429)  = ~\3926GAT(1420)  & ~\3742GAT(1328) ,
  \2507GAT(808)  = ~\843GAT(187)  & ~\2438GAT(776) ,
  \3944GAT(1403)  = ~\3894GAT(1367)  & ~\3893GAT(1366) ,
  \2221GAT(641)  = ~\2145GAT(623)  & ~\1272GAT(44) ,
  \1615GAT(411)  = ~\1567GAT(371)  & ~\1566GAT(370) ,
  \6220GAT(2413)  = \[23] ,
  \2523GAT(797)  = ~\2450GAT(773)  & ~\2305GAT(707) ,
  \1695GAT(460)  = ~\1528GAT(393)  & ~\1644GAT(435) ,
  \759GAT(215)  = \409GAT(24)  & \69GAT(4) ,
  \3500GAT(1246)  = ~\756GAT(216)  & ~\3433GAT(1212) ,
  \4302GAT(1592)  = ~\4185GAT(1546)  & ~\4248GAT(1567) ,
  \6014GAT(2322)  = ~\732GAT(224)  & ~\5981GAT(2304) ,
  \3338GAT(1167)  = ~\3177GAT(1090)  & ~\3292GAT(1141) ,
  \885GAT(173)  = \307GAT(18)  & \120GAT(7) ,
  \3408GAT(1178)  = ~\3356GAT(1152)  & ~\3314GAT(1132) ,
  \3591GAT(1268)  = ~\1143GAT(87)  & ~\3536GAT(1230) ,
  \1149GAT(85)  = \443GAT(26)  & \205GAT(12) ,
  \4178GAT(1536)  = ~\4114GAT(1515)  & ~\4055GAT(1490) ,
  \744GAT(220)  = \324GAT(19)  & \69GAT(4) ,
  \5804GAT(2225)  = ~\5749GAT(2204)  & ~\5752GAT(2203) ,
  \5844GAT(2251)  = ~\5792GAT(2235)  & ~\5740GAT(2206) ,
  \663GAT(247)  = \409GAT(24)  & \35GAT(2) ,
  \5639GAT(2147)  = ~\5569GAT(2131)  & ~\5395GAT(2045) ,
  \2745GAT(925)  = ~\558GAT(282)  & ~\2694GAT(906) ,
  \1143GAT(87)  = \409GAT(24)  & \205GAT(12) ,
  \1140GAT(88)  = \392GAT(23)  & \205GAT(12) ,
  \2661GAT(875)  = ~\2611GAT(854)  & ~\2561GAT(835) ,
  \3559GAT(1272)  = ~\3495GAT(1248)  & ~\3494GAT(1233) ,
  \2660GAT(884)  = ~\2493GAT(815)  & ~\2607GAT(855) ,
  \6026GAT(2315)  = ~\5990GAT(2302)  & ~\5993GAT(2301) ,
  \3521GAT(1234)  = ~\3449GAT(1208)  & ~\3296GAT(1140) ,
  \1137GAT(89)  = \375GAT(22)  & \205GAT(12) ,
  \5740GAT(2206)  = ~\5684GAT(2183)  & ~\5683GAT(2182) ,
  \1470GAT(356)  = ~\834GAT(190)  & ~\1419GAT(341) ,
  \2033GAT(580)  = ~\1224GAT(60)  & ~\2001GAT(562) ,
  \6281GAT(2442)  = ~\6277GAT(2439)  & ~\5727GAT(2167) ,
  \4571GAT(1687)  = ~\1056GAT(116)  & ~\4503GAT(1661) ,
  \2365GAT(762)  = ~\2329GAT(744)  & ~\2328GAT(740) ,
  \4711GAT(1774)  = ~\4531GAT(1698)  & ~\4650GAT(1746) ,
  \5401GAT(2042)  = ~\5344GAT(2018)  & ~\5343GAT(2017) ,
  \5009GAT(1901)  = ~\4886GAT(1851)  & ~\4950GAT(1873) ,
  \4622GAT(1709)  = ~\4566GAT(1689)  & ~\4380GAT(1602) ,
  \1886GAT(507)  = ~\1811GAT(488)  & ~\1676GAT(427) ,
  \4225GAT(1533)  = ~\1101GAT(101)  & ~\4155GAT(1508) ,
  \5213GAT(1961)  = ~\5151GAT(1950)  & ~\5094GAT(1910) ,
  \2826GAT(943)  = ~\2761GAT(921)  & ~\2706GAT(902) ,
  \3177GAT(1090)  = ~\3107GAT(1062)  & ~\2954GAT(995) ,
  \3095GAT(1065)  = ~\753GAT(217)  & ~\3040GAT(1046) ,
  \1783GAT(495)  = ~\789GAT(205)  & ~\1732GAT(478) ,
  \2344GAT(724)  = ~\2305GAT(707)  & ~\2251GAT(690) ,
  \1971GAT(571)  = ~\1856GAT(525)  & ~\1920GAT(554) ,
  \897GAT(169)  = \375GAT(22)  & \120GAT(7) ,
  \2822GAT(958)  = ~\702GAT(234)  & ~\2757GAT(922) ,
  \5599GAT(2111)  = ~\5536GAT(2102)  & ~\5535GAT(2086) ,
  \5817GAT(2221)  = ~\5764GAT(2209)  & ~\5706GAT(2174) ,
  \942GAT(154)  = \358GAT(21)  & \137GAT(8) ,
  \5323GAT(2025)  = ~\5194GAT(1967)  & ~\5262GAT(1992) ,
  \1851GAT(528)  = ~\1783GAT(495)  & ~\1648GAT(434) ,
  \2962GAT(993)  = ~\2853GAT(939)  & ~\2905GAT(971) ,
  \5650GAT(2144)  = ~\5516GAT(2092)  & ~\5581GAT(2117) ,
  \2224GAT(699)  = ~\2155GAT(681)  & ~\2154GAT(675) ,
  \4055GAT(1490)  = ~\4008GAT(1470)  & ~\4007GAT(1461) ,
  \2347GAT(727)  = ~\2201GAT(653)  & ~\2309GAT(706) ,
  \4061GAT(1488)  = ~\4012GAT(1468)  & ~\4011GAT(1459) ,
  \5451GAT(2068)  = ~\5333GAT(2021)  & ~\5395GAT(2045) ,
  \4973GAT(1877)  = ~\963GAT(147)  & ~\4916GAT(1844) ,
  \4595GAT(1720)  = ~\4535GAT(1697)  & ~\4534GAT(1685) ,
  \1696GAT(457)  = ~\1648GAT(434)  & ~\1597GAT(417) ,
  \4335GAT(1578)  = ~\4275GAT(1557)  & ~\4278GAT(1556) ,
  \3401GAT(1181)  = ~\3349GAT(1161)  & ~\3348GAT(1155) ,
  \4073GAT(1493)  = ~\906GAT(166)  & ~\4019GAT(1453) ,
  \6032GAT(2312)  = ~\6001GAT(2299)  & ~\6000GAT(2298) ,
  \5858GAT(2245)  = ~\5809GAT(2224)  & ~\5808GAT(2223) ,
  \747GAT(219)  = \341GAT(20)  & \69GAT(4) ,
  \2657GAT(879)  = ~\2603GAT(856)  & ~\2555GAT(837) ,
  \3111GAT(1061)  = ~\945GAT(153)  & ~\3052GAT(1040) ,
  \894GAT(170)  = \358GAT(21)  & \120GAT(7) ,
  \4384GAT(1600)  = ~\4335GAT(1578)  & ~\4278GAT(1556) ,
  \2142GAT(624)  = ~\2081GAT(609)  & ~\2080GAT(607) ,
  \1413GAT(343)  = ~\1380GAT(323)  & ~\1379GAT(324) ,
  \1885GAT(509)  = ~\1125GAT(93)  & ~\1811GAT(488) ,
  \3244GAT(1115)  = ~\3121GAT(1056)  & ~\3193GAT(1075) ,
  \5410GAT(2040)  = ~\5348GAT(2032)  & ~\5163GAT(1933) ,
  \4583GAT(1671)  = ~\4450GAT(1627)  & ~\4515GAT(1649) ,
  \2656GAT(886)  = ~\2483GAT(820)  & ~\2599GAT(857) ,
  \918GAT(162)  = \494GAT(29)  & \120GAT(7) ,
  \3612GAT(1293)  = ~\3491GAT(1249)  & ~\3559GAT(1272) ,
  \978GAT(142)  = \290GAT(17)  & \154GAT(9) ,
  \1920GAT(554)  = ~\1860GAT(524)  & ~\1859GAT(520) ,
  \5422GAT(2035)  = ~\5365GAT(2011)  & ~\5364GAT(2010) ,
  \1327GAT(298)  = ~\783GAT(207) ,
  \3055GAT(1039)  = ~\3006GAT(1017)  & ~\3005GAT(1010) ,
  \2700GAT(904)  = ~\2658GAT(885)  & ~\2657GAT(879) ,
  \2046GAT(619)  = ~\2011GAT(600)  & ~\2010GAT(597) ,
  \4461GAT(1624)  = ~\4350GAT(1573)  & ~\4401GAT(1595) ,
  \2030GAT(578)  = ~\2000GAT(564)  & ~\1999GAT(563) ,
  \4048GAT(1455)  = ~\1245GAT(53)  & ~\4001GAT(1433) ,
  \4554GAT(1680)  = ~\4487GAT(1662)  & ~\4486GAT(1659) ,
  \2823GAT(957)  = ~\2757GAT(922)  & ~\2607GAT(855) ,
  \4801GAT(1794)  = ~\1107GAT(99)  & ~\4742GAT(1767) ,
  \3494GAT(1233)  = ~\3429GAT(1213)  & ~\3374GAT(1191) ,
  \3533GAT(1221)  = ~\3466GAT(1200)  & ~\3465GAT(1199) ,
  \5825GAT(2218)  = ~\5770GAT(2197)  & ~\5773GAT(2196) ,
  \2635GAT(848)  = ~\2528GAT(794)  & ~\2579GAT(828) ,
  \3331GAT(1162)  = ~\3280GAT(1144)  & ~\3224GAT(1123) ,
  \5705GAT(2176)  = ~\5575GAT(2119)  & ~\5645GAT(2145) ,
  \4642GAT(1716)  = ~\1251GAT(51)  & ~\4587GAT(1682) ,
  \1053GAT(117)  = \443GAT(26)  & \171GAT(10) ,
  \5357GAT(2013)  = ~\5297GAT(1996)  & ~\5296GAT(1981) ,
  \5755GAT(2202)  = ~\5694GAT(2179)  & ~\5697GAT(2178) ,
  \1697GAT(458)  = ~\1533GAT(390)  & ~\1648GAT(434) ,
  \3830GAT(1385)  = ~\3764GAT(1364)  & ~\3709GAT(1341) ,
  \3049GAT(1041)  = ~\3002GAT(1021)  & ~\3001GAT(1012) ,
  \1600GAT(416)  = ~\1542GAT(386)  & ~\1541GAT(385) ,
  \1107GAT(99)  = \477GAT(28)  & \188GAT(11) ,
  \5831GAT(2215)  = ~\5781GAT(2194)  & ~\5780GAT(2193) ,
  \3923GAT(1410)  = ~\3873GAT(1374)  & ~\3872GAT(1373) ,
  \618GAT(262)  = \426GAT(25)  & \18GAT(1) ,
  \3361GAT(1151)  = ~\3254GAT(1111)  & ~\3317GAT(1131) ,
  \678GAT(242)  = \494GAT(29)  & \35GAT(2) ,
  \3221GAT(1124)  = ~\3161GAT(1100)  & ~\3160GAT(1085) ,
  \2712GAT(900)  = ~\2666GAT(878)  & ~\2665GAT(871) ,
  \5938GAT(2288)  = ~\5891GAT(2274)  & ~\5890GAT(2271) ,
  \2579GAT(828)  = ~\2532GAT(793)  & ~\2531GAT(788) ,
  \3902GAT(1419)  = ~\3841GAT(1396)  & ~\3840GAT(1383) ,
  \3505GAT(1244)  = ~\804GAT(200)  & ~\3437GAT(1211) ,
  \5214GAT(1971)  = ~\1014GAT(130)  & ~\5151GAT(1950) ,
  \3628GAT(1289)  = ~\3511GAT(1240)  & ~\3571GAT(1266) ,
  \4172GAT(1495)  = ~\4049GAT(1444)  & ~\4106GAT(1472) ,
  \3658GAT(1278)  = ~\3542GAT(1219)  & ~\3598GAT(1257) ,
  \5573GAT(2120)  = ~\5510GAT(2107)  & ~\5452GAT(2066) ,
  \4956GAT(1870)  = ~\4900GAT(1846)  & ~\4899GAT(1836) ,
  \828GAT(192)  = \528GAT(31)  & \86GAT(5) ,
  \3127GAT(1054)  = ~\3064GAT(1037)  & ~\3067GAT(1036) ,
  \4241GAT(1572)  = \[9] ,
  \888GAT(172)  = \324GAT(19)  & \120GAT(7) ,
  \4851GAT(1806)  = ~\4792GAT(1785)  & ~\4791GAT(1784) ,
  \3739GAT(1329)  = ~\3686GAT(1310)  & ~\3685GAT(1302) ,
  \4090GAT(1478)  = ~\3986GAT(1429)  & ~\4034GAT(1449) ,
  \2655GAT(881)  = ~\2599GAT(857)  & ~\2552GAT(838) ,
  \4737GAT(1755)  = ~\4683GAT(1732)  & ~\4625GAT(1708) ,
  \4566GAT(1689)  = ~\1008GAT(132)  & ~\4500GAT(1653) ,
  \2109GAT(634)  = ~\840GAT(188)  & ~\2055GAT(616) ,
  \3860GAT(1377)  = ~\3788GAT(1358)  & ~\3727GAT(1332) ,
  \2346GAT(722)  = ~\2309GAT(706)  & ~\2254GAT(689) ,
  \5898GAT(2268)  = ~\5846GAT(2250)  & ~\5849GAT(2249) ,
  \4604GAT(1715)  = ~\4550GAT(1691)  & ~\4549GAT(1681) ,
  \2289GAT(711)  = ~\2176GAT(668)  & ~\2239GAT(694) ,
  \660GAT(248)  = \392GAT(23)  & \35GAT(2) ,
  \1726GAT(480)  = ~\1693GAT(462)  & ~\1692GAT(461) ,
  \2251GAT(690)  = ~\2200GAT(655)  & ~\2199GAT(648) ,
  \3310GAT(1137)  = ~\1140GAT(88)  & ~\3248GAT(1121) ,
  \4793GAT(1783)  = ~\4738GAT(1756)  & ~\4737GAT(1755) ,
  \4290GAT(1564)  = ~\1248GAT(52)  & ~\4238GAT(1517) ,
  \1884GAT(505)  = ~\1811GAT(488)  & ~\1753GAT(471) ,
  \3368GAT(1194)  = ~\3326GAT(1175)  & ~\3325GAT(1168) ,
  \6225GAT(2415)  = ~\6221GAT(2412)  & ~\6002GAT(2297) ,
  \3842GAT(1395)  = ~\3772GAT(1362)  & ~\3616GAT(1292) ,
  \3747GAT(1327)  = ~\3647GAT(1281)  & ~\3693GAT(1299) ,
  \1095GAT(103)  = \409GAT(24)  & \188GAT(11) ,
  \3322GAT(1130)  = ~\3208GAT(1070)  & ~\3260GAT(1109) ,
  \4524GAT(1688)  = ~\4462GAT(1668)  & ~\4405GAT(1643) ,
  \6211GAT(2407)  = ~\6207GAT(2404)  & ~\6032GAT(2312) ,
  \3931GAT(1418)  = ~\1098GAT(102)  & ~\3877GAT(1382) ,
  \4357GAT(1612)  = ~\4302GAT(1592)  & ~\4248GAT(1567) ,
  \4173GAT(1537)  = ~\4110GAT(1516)  & ~\4052GAT(1491) ,
  \3699GAT(1296)  = ~\3658GAT(1278)  & ~\3657GAT(1277) ,
  \1987GAT(567)  = ~\1876GAT(513)  & ~\1932GAT(550) ,
  \5581GAT(2117)  = ~\5516GAT(2092)  & ~\5519GAT(2091) ,
  \3896GAT(1422)  = ~\3831GAT(1400)  & ~\3830GAT(1385) ,
  \1850GAT(530)  = ~\789GAT(205)  & ~\1783GAT(495) ,
  \2654GAT(887)  = ~\2478GAT(822)  & ~\2595GAT(858) ,
  \4578GAT(1672)  = ~\4509GAT(1651)  & ~\4512GAT(1650) ,
  \3712GAT(1339)  = ~\3667GAT(1320)  & ~\3666GAT(1311) ,
  \4689GAT(1729)  = ~\4633GAT(1706)  & ~\4632GAT(1705) ,
  \5230GAT(1970)  = ~\1209GAT(65)  & ~\5169GAT(1930) ,
  \5032GAT(1890)  = ~\4968GAT(1878)  & ~\4787GAT(1786) ,
  \2706GAT(902)  = ~\2662GAT(882)  & ~\2661GAT(875) ,
  \708GAT(232)  = \392GAT(23)  & \52GAT(3) ,
  \1698GAT(455)  = ~\1652GAT(433)  & ~\1600GAT(416) ,
  \1407GAT(345)  = ~\1376GAT(327)  & ~\1375GAT(328) ,
  \2650GAT(841)  = ~\2591GAT(829)  & ~\2410GAT(746) ,
  \4237GAT(1519)  = ~\4100GAT(1474)  & ~\4167GAT(1496) ,
  \3562GAT(1271)  = ~\3500GAT(1246)  & ~\3499GAT(1232) ,
  \2518GAT(800)  = ~\2446GAT(774)  & ~\2301GAT(708) ,
  \3157GAT(1101)  = ~\3091GAT(1066)  & ~\2938GAT(999) ,
  \4058GAT(1489)  = ~\4010GAT(1469)  & ~\4009GAT(1460) ,
  \2999GAT(1014)  = ~\2950GAT(996)  & ~\2896GAT(976) ,
  \3193GAT(1075)  = ~\3121GAT(1056)  & ~\3124GAT(1055) ,
  \756GAT(216)  = \392GAT(23)  & \69GAT(4) ,
  \2227GAT(698)  = ~\2160GAT(679)  & ~\2159GAT(672) ,
  \1029GAT(125)  = \307GAT(18)  & \171GAT(10) ,
  \4456GAT(1625)  = ~\4395GAT(1597)  & ~\4398GAT(1596) ,
  \3280GAT(1144)  = ~\3162GAT(1099)  & ~\3224GAT(1123) ,
  \1664GAT(430)  = ~\1553GAT(378)  & ~\1609GAT(413) ,
  \1089GAT(105)  = \375GAT(22)  & \188GAT(11) ,
  \2539GAT(786)  = ~\2464GAT(768)  & ~\2467GAT(767) ,
  \3821GAT(1344)  = ~\3757GAT(1323)  & ~\1290GAT(38) ,
  \3813GAT(1347)  = ~\3751GAT(1335)  & ~\3699GAT(1296) ,
  \2878GAT(982)  = ~\2812GAT(962)  & ~\2811GAT(952) ,
  \4220GAT(1535)  = ~\1053GAT(117)  & ~\4152GAT(1500) ,
  \1699GAT(456)  = ~\1538GAT(387)  & ~\1652GAT(433) ,
  \4414GAT(1638)  = ~\4360GAT(1619)  & ~\4359GAT(1610) ,
  \2166GAT(674)  = ~\2097GAT(637)  & ~\1959GAT(574) ,
  \585GAT(273)  = \511GAT(30)  & \1GAT(0) ,
  \1410GAT(344)  = ~\1378GAT(325)  & ~\1377GAT(326) ,
  \3004GAT(1019)  = ~\2848GAT(942)  & ~\2958GAT(994) ,
  \4932GAT(1825)  = ~\4866GAT(1802)  & ~\4805GAT(1780) ,
  \2392GAT(751)  = ~\2347GAT(727)  & ~\2346GAT(722) ,
  \2164GAT(669)  = ~\2097GAT(637)  & ~\2046GAT(619) ,
  \4031GAT(1450)  = ~\3985GAT(1434)  & ~\3984GAT(1430) ,
  \2434GAT(777)  = ~\795GAT(203)  & ~\2377GAT(758) ,
  \975GAT(143)  = \273GAT(16)  & \154GAT(9) ,
  \4802GAT(1781)  = ~\4742GAT(1767)  & ~\4578GAT(1672) ,
  \6286GAT(2446)  = ~\6277GAT(2439)  & ~\6281GAT(2442) ,
  \2149GAT(678)  = ~\2085GAT(640)  & ~\2037GAT(622) ,
  \5941GAT(2287)  = ~\5892GAT(2270)  & ~\5895GAT(2269) ,
  \3233GAT(1118)  = ~\3181GAT(1089)  & ~\3180GAT(1079) ,
  \1923GAT(553)  = ~\1865GAT(521)  & ~\1864GAT(517) ,
  \4833GAT(1817)  = ~\768GAT(212)  & ~\4772GAT(1790) ,
  \5409GAT(2051)  = ~\1113GAT(97)  & ~\5348GAT(2032) ,
  \4964GAT(1868)  = ~\4839GAT(1811)  & ~\4907GAT(1834) ,
  \3404GAT(1180)  = ~\3350GAT(1154)  & ~\3353GAT(1153) ,
  \4078GAT(1492)  = ~\954GAT(150)  & ~\4022GAT(1464) ,
  \3334GAT(1171)  = ~\3167GAT(1096)  & ~\3284GAT(1143) ,
  \5866GAT(2254)  = ~\972GAT(144)  & ~\5813GAT(2233) ,
  \5184GAT(1975)  = ~\675GAT(243)  & ~\5124GAT(1946) ,
  \2368GAT(761)  = ~\2331GAT(743)  & ~\2330GAT(738) ,
  \6231GAT(2417)  = ~\6227GAT(2414)  & ~\5968GAT(2277) ,
  \5092GAT(1911)  = ~\5038GAT(1888)  & ~\4977GAT(1863) ,
  \3070GAT(1035)  = ~\3016GAT(1007)  & ~\3019GAT(1006) ,
  \6102GAT(2349)  = ~\6046GAT(2330)  & ~\6076GAT(2340) ,
  \4858GAT(1805)  = ~\4796GAT(1796)  & ~\4739GAT(1754) ,
  \6002GAT(2297)  = ~\5967GAT(2279)  & ~\5966GAT(2278) ,
  \3180GAT(1079)  = ~\3111GAT(1061)  & ~\3052GAT(1040) ,
  \6124GAT(2367)  = ~\6108GAT(2362)  & ~\6111GAT(2360) ,
  \5073GAT(1917)  = ~\5022GAT(1898)  & ~\5021GAT(1893) ,
  \6090GAT(2354)  = ~\636GAT(256)  & ~\6064GAT(2346) ,
  \4507GAT(1652)  = ~\4444GAT(1641)  & ~\4386GAT(1599) ,
  \2990GAT(1030)  = ~\2813GAT(961)  & ~\2930GAT(1001) ,
  \2757GAT(922)  = ~\702GAT(234)  & ~\2703GAT(903) ,
  \6040GAT(2335)  = ~\684GAT(240)  & ~\6011GAT(2319) ,
  \3062GAT(1038)  = ~\3010GAT(1015)  & ~\2968GAT(988) ,
  \675GAT(243)  = \477GAT(28)  & \35GAT(2) ,
  \2831GAT(940)  = ~\2765GAT(920)  & ~\2709GAT(901) ,
  \5933GAT(2289)  = ~\5886GAT(2275)  & ~\5837GAT(2252) ,
  \5683GAT(2182)  = ~\5624GAT(2152)  & ~\5557GAT(2125) ,
  \1811GAT(488)  = ~\1125GAT(93)  & ~\1753GAT(471) ,
  \5226GAT(1957)  = ~\5103GAT(1908)  & ~\5163GAT(1933) ,
  \4899GAT(1836)  = ~\4833GAT(1817)  & ~\4772GAT(1790) ,
  \6207GAT(2404)  = ~\6201GAT(2402)  & ~\5996GAT(2300) ,
  \4854GAT(1815)  = ~\1011GAT(131)  & ~\4793GAT(1783) ,
  \1323GAT(299)  = ~\735GAT(223) ,
  \4327GAT(1581)  = ~\4269GAT(1571)  & ~\4217GAT(1524) ,
  \3040GAT(1046)  = ~\2996GAT(1027)  & ~\2995GAT(1018) ,
  \3653GAT(1279)  = ~\3592GAT(1259)  & ~\3595GAT(1258) ,
  \3942GAT(1404)  = ~\3889GAT(1368)  & ~\3818GAT(1345) ,
  \6130GAT(2364)  = ~\6119GAT(2358)  & ~\6118GAT(2357) ,
  \3224GAT(1123)  = ~\3166GAT(1098)  & ~\3165GAT(1083) ,
  \900GAT(168)  = \392GAT(23)  & \120GAT(7) ,
  \1603GAT(415)  = ~\1547GAT(383)  & ~\1546GAT(382) ,
  \3141GAT(1108)  = ~\561GAT(281)  & ~\3079GAT(1069) ,
  \4232GAT(1520)  = ~\4161GAT(1498)  & ~\4164GAT(1497) ,
  \732GAT(224)  = \528GAT(31)  & \52GAT(3) ,
  \3254GAT(1111)  = ~\3202GAT(1080)  & ~\3022GAT(1005) ,
  \3260GAT(1109)  = ~\3208GAT(1070)  & ~\1284GAT(40) ,
  \4953GAT(1871)  = ~\4895GAT(1848)  & ~\4894GAT(1838) ,
  \1779GAT(496)  = ~\741GAT(221)  & ~\1729GAT(479) ,
  \5467GAT(2062)  = ~\5410GAT(2040)  & ~\5413GAT(2039) ,
  \1404GAT(346)  = ~\1374GAT(329)  & ~\1373GAT(330) ,
  \4007GAT(1461)  = ~\3951GAT(1442)  & ~\3899GAT(1421) ,
  \4106GAT(1472)  = ~\4049GAT(1444)  & ~\1293GAT(37) ,
  \1889GAT(503)  = ~\1815GAT(487)  & ~\1756GAT(469) ,
  \4411GAT(1640)  = ~\4358GAT(1620)  & ~\4357GAT(1612) ,
  \6069GAT(2345)  = ~\684GAT(240)  & ~\6040GAT(2335) ,
  \2977GAT(986)  = ~\2917GAT(974)  & ~\2739GAT(890) ,
  \1648GAT(434)  = ~\1533GAT(390)  & ~\1597GAT(417) ,
  \2744GAT(889)  = ~\2650GAT(841)  & ~\2690GAT(859) ,
  \2837GAT(950)  = ~\846GAT(186)  & ~\2769GAT(919) ,
  \1652GAT(433)  = ~\1538GAT(387)  & ~\1600GAT(416) ,
  \2422GAT(780)  = ~\651GAT(251)  & ~\2368GAT(761) ,
  \4717GAT(1771)  = ~\4546GAT(1692)  & ~\4662GAT(1743) ,
  \3845GAT(1381)  = ~\3776GAT(1361)  & ~\3718GAT(1337) ,
  \2064GAT(613)  = ~\2023GAT(588)  & ~\2022GAT(585) ,
  \5972GAT(2308)  = ~\5934GAT(2294)  & ~\5933GAT(2289) ,
  \5327GAT(2034)  = ~\870GAT(178)  & ~\5268GAT(1989) ,
  \4423GAT(1645)  = ~\861GAT(181)  & ~\4365GAT(1606) ,
  \5455GAT(2079)  = ~\1017GAT(129)  & ~\5401GAT(2042) ,
  \5005GAT(1902)  = ~\4881GAT(1853)  & ~\4947GAT(1875) ,
  \2508GAT(806)  = ~\2438GAT(776)  & ~\2293GAT(710) ,
  \2165GAT(676)  = ~\696GAT(236)  & ~\2097GAT(637) ,
  \6261GAT(2432)  = ~\6257GAT(2429)  & ~\5831GAT(2215) ,
  \5553GAT(2132)  = ~\726GAT(226)  & ~\5489GAT(2109) ,
  \4779GAT(1789)  = ~\4721GAT(1770)  & ~\4668GAT(1736) ,
  \3392GAT(1192)  = ~\996GAT(136)  & ~\3341GAT(1156) ,
  \903GAT(167)  = \409GAT(24)  & \120GAT(7) ,
  \3389GAT(1184)  = ~\3340GAT(1165)  & ~\3339GAT(1157) ,
  \3797GAT(1352)  = ~\3735GAT(1340)  & ~\3734GAT(1331) ,
  \2761GAT(921)  = ~\750GAT(218)  & ~\2706GAT(902) ,
  \2105GAT(635)  = ~\792GAT(204)  & ~\2052GAT(617) ,
  \3664GAT(1313)  = ~\3608GAT(1294)  & ~\3556GAT(1273) ,
  \5389GAT(2047)  = ~\5327GAT(2034)  & ~\5142GAT(1940) ,
  \3735GAT(1340)  = ~\999GAT(135)  & ~\3681GAT(1312) ,
  \3003GAT(1011)  = ~\2958GAT(994)  & ~\2902GAT(973) ,
  \3007GAT(1009)  = ~\2967GAT(992)  & ~\2966GAT(989) ,
  \1839GAT(532)  = ~\1775GAT(497)  & ~\1726GAT(480) ,
  \5595GAT(2128)  = ~\1212GAT(64)  & ~\5531GAT(2104) ,
  \3727GAT(1332)  = ~\3677GAT(1314)  & ~\3676GAT(1304) ,
  \3757GAT(1323)  = ~\3702GAT(1305)  & ~\3548GAT(1217) ,
  \2576GAT(830)  = ~\2527GAT(796)  & ~\2526GAT(789) ,
  \1486GAT(352)  = ~\1026GAT(126)  & ~\1431GAT(337) ,
  \1836GAT(537)  = ~\1771GAT(498)  & ~\1636GAT(437) ,
  \5043GAT(1887)  = ~\4922GAT(1829)  & ~\4980GAT(1862) ,
  \6236GAT(2421)  = ~\6227GAT(2414)  & ~\6231GAT(2417) ,
  \3099GAT(1064)  = ~\801GAT(201)  & ~\3043GAT(1044) ,
  \3670GAT(1308)  = ~\3620GAT(1291)  & ~\3565GAT(1269) ,
  \3323GAT(1170)  = ~\3264GAT(1148)  & ~\3212GAT(1127) ,
  \4775GAT(1798)  = ~\816GAT(196)  & ~\4718GAT(1761) ,
  \4563GAT(1676)  = ~\4499GAT(1655)  & ~\4498GAT(1654) ,
  \5056GAT(1882)  = ~\4994GAT(1872)  & ~\4993GAT(1858) ,
  \588GAT(272)  = \528GAT(31)  & \1GAT(0) ,
  \2285GAT(712)  = ~\2171GAT(671)  & ~\2236GAT(695) ,
  \1807GAT(489)  = ~\1077GAT(109)  & ~\1750GAT(472) ,
  \4028GAT(1451)  = ~\3980GAT(1435)  & ~\3800GAT(1351) ,
  \2627GAT(850)  = ~\2518GAT(800)  & ~\2573GAT(831) ,
  \2659GAT(877)  = ~\2607GAT(855)  & ~\2558GAT(836) ,
  \5780GAT(2193)  = ~\5721GAT(2170)  & ~\5663GAT(2139) ,
  \4339GAT(1576)  = ~\4281GAT(1555)  & ~\4229GAT(1521) ,
  \3602GAT(1255)  = ~\3548GAT(1217)  & ~\1287GAT(39) ,
  \3198GAT(1074)  = ~\3064GAT(1037)  & ~\3127GAT(1054) ,
  \825GAT(193)  = \511GAT(30)  & \86GAT(5) ,
  \4541GAT(1694)  = ~\4474GAT(1665)  & ~\4306GAT(1591) ,
  \4217GAT(1524)  = ~\4151GAT(1502)  & ~\4150GAT(1501) ,
  \2169GAT(666)  = ~\2101GAT(636)  & ~\2049GAT(618) ,
  \2313GAT(705)  = ~\2206GAT(650)  & ~\2257GAT(688) ,
  \5968GAT(2277)  = ~\5924GAT(2260)  & ~\5923GAT(2259) ,
  \4194GAT(1543)  = ~\762GAT(214)  & ~\4126GAT(1512) ,
  \3702GAT(1305)  = ~\1242GAT(54)  & ~\3659GAT(1276) ,
  \3911GAT(1415)  = ~\3856GAT(1390)  & ~\3855GAT(1378) ,
  \3353GAT(1153)  = ~\3310GAT(1137)  & ~\3309GAT(1134) ,
  \3115GAT(1060)  = ~\993GAT(137)  & ~\3055GAT(1039) ,
  \3852GAT(1391)  = ~\3780GAT(1360)  & ~\3624GAT(1290) ,
  \6160GAT(2383)  = \[17] ,
  \5787GAT(2230)  = ~\5734GAT(2213)  & ~\5676GAT(2185) ,
  \3236GAT(1117)  = ~\3186GAT(1086)  & ~\3185GAT(1077) ,
  \2658GAT(885)  = ~\2488GAT(818)  & ~\2603GAT(856) ,
  \4725GAT(1760)  = ~\4671GAT(1741)  & ~\4613GAT(1711) ,
  \4140GAT(1505)  = ~\4073GAT(1493)  & ~\3917GAT(1413) ,
  \3894GAT(1367)  = ~\3757GAT(1323)  & ~\3821GAT(1344) ,
  \855GAT(183)  = \409GAT(24)  & \103GAT(6) ,
  \981GAT(141)  = \307GAT(18)  & \154GAT(9) ,
  \4758GAT(1748)  = ~\4704GAT(1725)  & ~\1299GAT(35) ,
  \2975GAT(987)  = ~\2917GAT(974)  & ~\2870GAT(926) ,
  \5064GAT(1880)  = ~\4943GAT(1822)  & ~\5001GAT(1855) ,
  \1098GAT(102)  = \426GAT(25)  & \188GAT(11) ,
  \4453GAT(1626)  = ~\4394GAT(1609)  & ~\4393GAT(1598) ,
  \4362GAT(1618)  = ~\4195GAT(1542)  & ~\4310GAT(1590) ,
  \2709GAT(901)  = ~\2664GAT(880)  & ~\2663GAT(873) ,
  \5365GAT(2011)  = ~\5236GAT(1953)  & ~\5304GAT(1978) ,
  \4229GAT(1521)  = ~\4160GAT(1507)  & ~\4159GAT(1499) ,
  \1729GAT(479)  = ~\1695GAT(460)  & ~\1694GAT(459) ,
  \2438GAT(776)  = ~\843GAT(187)  & ~\2380GAT(757) ,
  \1059GAT(115)  = \477GAT(28)  & \171GAT(10) ,
  \4814GAT(1776)  = ~\4759GAT(1749)  & ~\4758GAT(1748) ,
  \5106GAT(1907)  = ~\5052GAT(1894)  & ~\5051GAT(1884) ,
  \882GAT(174)  = \290GAT(17)  & \120GAT(7) ,
  \5315GAT(2027)  = ~\5255GAT(2003)  & ~\5254GAT(1994) ,
  \4912GAT(1833)  = ~\4781GAT(1788)  & ~\4845GAT(1809) ,
  \4500GAT(1653)  = ~\4440GAT(1631)  & ~\4439GAT(1630) ,
  \705GAT(233)  = \375GAT(22)  & \52GAT(3) ,
  \5633GAT(2160)  = ~\873GAT(177)  & ~\5566GAT(2121) ,
  \3581GAT(1262)  = ~\3527GAT(1224)  & ~\3458GAT(1202) ,
  \3160GAT(1085)  = ~\3095GAT(1065)  & ~\3040GAT(1046) ,
  \2478GAT(822)  = ~\2414GAT(782)  & ~\2269GAT(716) ,
  \2532GAT(793)  = ~\1083GAT(107)  & ~\2458GAT(771) ,
  \2921GAT(966)  = ~\2873GAT(932)  & ~\2803GAT(907) ,
  \2170GAT(673)  = ~\744GAT(220)  & ~\2101GAT(636) ,
  \2374GAT(759)  = ~\2335GAT(739)  & ~\2334GAT(734) ,
  \2549GAT(839)  = ~\2482GAT(821)  & ~\2481GAT(813) ,
  \3636GAT(1284)  = ~\3577GAT(1264)  & ~\3524GAT(1225) ,
  \6097GAT(2350)  = ~\6070GAT(2342)  & ~\6073GAT(2341) ,
  \4251GAT(1566)  = ~\4194GAT(1543)  & ~\4193GAT(1531) ,
  \3989GAT(1428)  = ~\3931GAT(1418)  & ~\3930GAT(1409) ,
  \5151GAT(1950)  = ~\1014GAT(130)  & ~\5094GAT(1910) ,
  \6035GAT(2333)  = ~\6005GAT(2324)  & ~\5972GAT(2308) ,
  \5979GAT(2305)  = ~\5941GAT(2287)  & ~\5895GAT(2269) ,
  \4821GAT(1820)  = ~\624GAT(260)  & ~\4763GAT(1793) ,
  \4344GAT(1585)  = ~\1200GAT(68)  & ~\4287GAT(1552) ,
  \2533GAT(791)  = ~\2458GAT(771)  & ~\2313GAT(705) ,
  \1859GAT(520)  = ~\1791GAT(493)  & ~\1738GAT(476) ,
  \6019GAT(2321)  = ~\780GAT(208)  & ~\5984GAT(2311) ,
  \6057GAT(2327)  = ~\5990GAT(2302)  & ~\6026GAT(2315) ,
  \2548GAT(840)  = \[4] ,
  \2171GAT(671)  = ~\2101GAT(636)  & ~\1963GAT(573) ,
  \4089GAT(1477)  = ~\4034GAT(1449)  & ~\3989GAT(1428) ,
  \2922GAT(972)  = ~\1233GAT(57)  & ~\2873GAT(932) ,
  \6180GAT(2393)  = \[19] ,
  \2067GAT(612)  = ~\2025GAT(586)  & ~\2024GAT(583) ,
  \4920GAT(1830)  = ~\4854GAT(1815)  & ~\4793GAT(1783) ,
  \1834GAT(535)  = ~\1771GAT(498)  & ~\1723GAT(481) ,
  \3172GAT(1093)  = ~\3103GAT(1063)  & ~\2950GAT(996) ,
  \5383GAT(2054)  = ~\822GAT(194)  & ~\5324GAT(2023) ,
  \3151GAT(1104)  = ~\657GAT(249)  & ~\3087GAT(1067) ,
  \993GAT(137)  = \375GAT(22)  & \154GAT(9) ,
  \4155GAT(1508)  = ~\1101GAT(101)  & ~\4091GAT(1476) ,
  \1835GAT(539)  = ~\645GAT(253)  & ~\1771GAT(498) ,
  \5380GAT(2049)  = ~\5323GAT(2025)  & ~\5322GAT(2024) ,
  \783GAT(207)  = \273GAT(16)  & \86GAT(5) ,
  \1775GAT(497)  = ~\693GAT(237)  & ~\1726GAT(480) ,
  \2001GAT(562)  = ~\1946GAT(546)  & ~\1945GAT(545) ,
  \4784GAT(1787)  = ~\4726GAT(1769)  & ~\4725GAT(1760) ,
  \3980GAT(1435)  = ~\1002GAT(134)  & ~\3923GAT(1410) ,
  \4643GAT(1702)  = ~\4587GAT(1682)  & ~\4401GAT(1595) ,
  \1644GAT(435)  = ~\1528GAT(393)  & ~\1594GAT(418) ,
  \5796GAT(2228)  = ~\5743GAT(2211)  & ~\5685GAT(2181) ,
  \4285GAT(1553)  = ~\4232GAT(1520)  & ~\4164GAT(1497) ,
  \4968GAT(1878)  = ~\915GAT(163)  & ~\4913GAT(1831) ,
  \4011GAT(1459)  = ~\3959GAT(1440)  & ~\3905GAT(1417) ,
  \3197GAT(1073)  = ~\3127GAT(1054)  & ~\3067GAT(1036) ,
  \2145GAT(623)  = ~\2082GAT(606)  & ~\1272GAT(44) ,
  \3831GAT(1400)  = ~\615GAT(263)  & ~\3764GAT(1364) ,
  \3685GAT(1302)  = ~\3641GAT(1286)  & ~\3583GAT(1261) ,
  \3326GAT(1175)  = ~\3147GAT(1105)  & ~\3268GAT(1147) ,
  \1026GAT(126)  = \290GAT(17)  & \171GAT(10) ,
  \693GAT(237)  = \307GAT(18)  & \52GAT(3) ,
  \669GAT(245)  = \443GAT(26)  & \35GAT(2) ,
  \3272GAT(1146)  = ~\3152GAT(1103)  & ~\3218GAT(1125) ,
  \5564GAT(2122)  = ~\5501GAT(2097)  & ~\5443GAT(2070) ,
  \990GAT(138)  = \358GAT(21)  & \154GAT(9) ,
  \4536GAT(1696)  = ~\4470GAT(1666)  & ~\4302GAT(1592) ,
  \4361GAT(1608)  = ~\4310GAT(1590)  & ~\4254GAT(1565) ,
  \5053GAT(1883)  = ~\4989GAT(1874)  & ~\4808GAT(1779) ,
  \4712GAT(1764)  = ~\4654GAT(1745)  & ~\4598GAT(1719) ,
  \4666GAT(1737)  = ~\4607GAT(1714)  & ~\4554GAT(1680) ,
  \5339GAT(2019)  = ~\5277GAT(1987)  & ~\5280GAT(1986) ,
  \6266GAT(2436)  = ~\6257GAT(2429)  & ~\6261GAT(2432) ,
  \2000GAT(564)  = ~\1891GAT(504)  & ~\1941GAT(547) ,
  \1419GAT(341)  = ~\1384GAT(319)  & ~\1383GAT(320) ,
  \3441GAT(1210)  = ~\852GAT(184)  & ~\3383GAT(1187) ,
  \6191GAT(2397)  = ~\6187GAT(2394)  & ~\6082GAT(2337) ,
  \3514GAT(1227)  = ~\3445GAT(1209)  & ~\3386GAT(1186) ,
  \2684GAT(861)  = ~\2644GAT(846)  & ~\2470GAT(766) ,
  \3074GAT(1033)  = ~\3022GAT(1005)  & ~\2980GAT(985) ,
  \2923GAT(965)  = ~\2873GAT(932)  & ~\2690GAT(859) ,
  \912GAT(164)  = \460GAT(27)  & \120GAT(7) ,
  \690GAT(238)  = \290GAT(17)  & \52GAT(3) ,
  \5176GAT(1977)  = ~\579GAT(275)  & ~\5118GAT(1948) ,
  \3356GAT(1152)  = ~\3311GAT(1133)  & ~\3314GAT(1132) ,
  \3772GAT(1362)  = ~\711GAT(231)  & ~\3715GAT(1338) ,
  \1632GAT(438)  = ~\1513GAT(402)  & ~\1585GAT(421) ,
  \5697GAT(2178)  = ~\5638GAT(2159)  & ~\5637GAT(2148) ,
  \5628GAT(2150)  = ~\5560GAT(2124)  & ~\5498GAT(2098) ,
  \5352GAT(2015)  = ~\5292GAT(1998)  & ~\5227GAT(1955) ,
  \6167GAT(2384)  = ~\6161GAT(2382)  & ~\6097GAT(2350) ,
  \2052GAT(617)  = ~\2015GAT(596)  & ~\2014GAT(593) ,
  \4697GAT(1738)  = ~\1203GAT(67)  & ~\4637GAT(1718) ,
  \1691GAT(464)  = ~\1518GAT(399)  & ~\1636GAT(437) ,
  \5913GAT(2263)  = ~\5861GAT(2255)  & ~\5700GAT(2177) ,
  \1609GAT(413)  = ~\1557GAT(377)  & ~\1556GAT(376) ,
  \2317GAT(702)  = ~\2260GAT(687)  & ~\2214GAT(644) ,
  \5296GAT(1981)  = ~\5230GAT(1970)  & ~\5169GAT(1930) ,
  \2377GAT(758)  = ~\2337GAT(737)  & ~\2336GAT(732) ,
  \2531GAT(788)  = ~\2458GAT(771)  & ~\2395GAT(750) ,
  \3540GAT(1220)  = ~\3470GAT(1206)  & ~\3410GAT(1177) ,
  \3465GAT(1199)  = ~\3404GAT(1180)  & ~\3353GAT(1153) ,
  \3340GAT(1165)  = ~\3182GAT(1087)  & ~\3296GAT(1140) ,
  \3748GAT(1325)  = ~\3698GAT(1298)  & ~\3697GAT(1297) ,
  \4319GAT(1588)  = ~\4205GAT(1538)  & ~\4260GAT(1562) ,
  \5180GAT(1976)  = ~\627GAT(259)  & ~\5121GAT(1947) ,
  \5277GAT(1987)  = ~\5209GAT(1972)  & ~\5038GAT(1888) ,
  \4474GAT(1665)  = ~\717GAT(229)  & ~\4414GAT(1638) ,
  \612GAT(264)  = \392GAT(23)  & \18GAT(1) ,
  \738GAT(222)  = \290GAT(17)  & \69GAT(4) ,
  \3930GAT(1409)  = ~\3877GAT(1382)  & ~\3806GAT(1348) ,
  \4813GAT(1778)  = ~\4698GAT(1727)  & ~\4754GAT(1750) ,
  \[0]  = \273GAT(16)  & \1GAT(0) ,
  \3825GAT(1387)  = ~\3760GAT(1365)  & ~\3706GAT(1343) ,
  \5654GAT(2158)  = ~\1116GAT(96)  & ~\5587GAT(2114) ,
  \[1]  = ~\1507GAT(407)  & ~\1506GAT(406) ,
  \3873GAT(1374)  = ~\3736GAT(1330)  & ~\3800GAT(1351) ,
  \5980GAT(2306)  = ~\5892GAT(2270)  & ~\5941GAT(2287) ,
  \4551GAT(1690)  = ~\4482GAT(1663)  & ~\4314GAT(1589) ,
  \2687GAT(860)  = ~\2649GAT(845)  & ~\2648GAT(842) ,
  \[2]  = ~\1825GAT(544)  & ~\1824GAT(541) ,
  \5413GAT(2039)  = ~\5353GAT(2030)  & ~\5352GAT(2015) ,
  \[3]  = ~\2150GAT(683)  & ~\2149GAT(678) ,
  \3780GAT(1360)  = ~\807GAT(199)  & ~\3721GAT(1336) ,
  \6155GAT(2380)  = ~\6151GAT(2377)  & ~\6135GAT(2369) ,
  \[4]  = ~\2477GAT(823)  & ~\2476GAT(816) ,
  \3855GAT(1378)  = ~\3784GAT(1359)  & ~\3724GAT(1334) ,
  \822GAT(194)  = \494GAT(29)  & \86GAT(5) ,
  \[5]  = ~\2807GAT(964)  & ~\2806GAT(955) ,
  \2938GAT(999)  = ~\2823GAT(957)  & ~\2887GAT(979) ,
  \5679GAT(2184)  = ~\5618GAT(2161)  & ~\5621GAT(2153) ,
  \[6]  = ~\3141GAT(1108)  & ~\3140GAT(1097) ,
  \3230GAT(1120)  = ~\3176GAT(1092)  & ~\3175GAT(1081) ,
  \2976GAT(990)  = ~\1185GAT(73)  & ~\2917GAT(974) ,
  \3317GAT(1131)  = ~\3254GAT(1111)  & ~\3257GAT(1110) ,
  \[7]  = ~\3480GAT(1254)  & ~\3479GAT(1241) ,
  \3484GAT(1238)  = ~\3421GAT(1215)  & ~\3368GAT(1194) ,
  \5425GAT(2077)  = ~\5366GAT(2058)  & ~\5309GAT(2029) ,
  \[8]  = ~\3826GAT(1402)  & ~\3825GAT(1387) ,
  \4746GAT(1753)  = ~\4692GAT(1739)  & ~\4634GAT(1704) ,
  \4016GAT(1466)  = ~\3852GAT(1391)  & ~\3967GAT(1438) ,
  \[9]  = ~\4174GAT(1551)  & ~\4173GAT(1537) ,
  \4150GAT(1501)  = ~\4085GAT(1479)  & ~\4031GAT(1450) ,
  \2989GAT(1024)  = ~\2930GAT(1001)  & ~\2881GAT(981) ,
  \720GAT(228)  = \460GAT(27)  & \52GAT(3) ,
  \2402GAT(749)  = ~\2353GAT(723)  & ~\2319GAT(701) ,
  \3016GAT(1007)  = ~\2971GAT(991)  & ~\2797GAT(910) ,
  \3662GAT(1315)  = ~\3604GAT(1295)  & ~\3553GAT(1274) ,
  \1690GAT(463)  = ~\1636GAT(437)  & ~\1588GAT(420) ,
  \780GAT(208)  = \528GAT(31)  & \69GAT(4) ,
  \1528GAT(393)  = ~\1462GAT(358)  & ~\1327GAT(298) ,
  \5155GAT(1936)  = ~\5097GAT(1923)  & ~\5044GAT(1885) ,
  \3300GAT(1136)  = ~\3239GAT(1116)  & ~\3190GAT(1076) ,
  \3947GAT(1443)  = ~\3827GAT(1401)  & ~\3896GAT(1422) ,
  \4870GAT(1800)  = ~\4808GAT(1779)  & ~\4751GAT(1751) ,
  \1855GAT(527)  = ~\837GAT(189)  & ~\1787GAT(494) ,
  \5204GAT(1963)  = ~\5142GAT(1940)  & ~\5085GAT(1914) ,
  \1056GAT(116)  = \460GAT(27)  & \171GAT(10) ,
  \2476GAT(816)  = ~\2414GAT(782)  & ~\2362GAT(763) ,
  \5167GAT(1931)  = ~\5109GAT(1906)  & ~\5056GAT(1882) ,
  \5097GAT(1923)  = ~\1062GAT(114)  & ~\5044GAT(1885) ,
  \666GAT(246)  = \426GAT(25)  & \35GAT(2) ,
  \5956GAT(2282)  = ~\5907GAT(2273)  & ~\5755GAT(2202) ,
  \5388GAT(2053)  = ~\870GAT(178)  & ~\5327GAT(2034) ,
  \3881GAT(1371)  = ~\3809GAT(1356)  & ~\3748GAT(1325) ,
  \1840GAT(536)  = ~\693GAT(237)  & ~\1775GAT(497) ,
  \5239GAT(1999)  = ~\5176GAT(1977)  & ~\5118GAT(1948) ,
  \5671GAT(2137)  = ~\5537GAT(2085)  & ~\5602GAT(2110) ,
  \924GAT(160)  = \528GAT(31)  & \120GAT(7) ,
  \5066GAT(1929)  = ~\4881GAT(1853)  & ~\5005GAT(1902) ,
  \2653GAT(883)  = ~\2595GAT(858)  & ~\2549GAT(839) ,
  \858GAT(182)  = \426GAT(25)  & \103GAT(6) ,
  \2994GAT(1028)  = ~\2823GAT(957)  & ~\2938GAT(999) ,
  \2887GAT(979)  = ~\2827GAT(956)  & ~\2826GAT(943) ,
  \3899GAT(1421)  = ~\3836GAT(1398)  & ~\3835GAT(1384) ,
  \6020GAT(2317)  = ~\5984GAT(2311)  & ~\5852GAT(2248) ,
  \582GAT(274)  = \494GAT(29)  & \1GAT(0) ,
  \6187GAT(2394)  = ~\6181GAT(2392)  & ~\6052GAT(2328) ,
  \3837GAT(1397)  = ~\3768GAT(1363)  & ~\3612GAT(1293) ,
  \5459GAT(2065)  = ~\5404GAT(2052)  & ~\5345GAT(2016) ,
  \3977GAT(1431)  = ~\3922GAT(1412)  & ~\3921GAT(1411) ,
  \2506GAT(798)  = ~\2438GAT(776)  & ~\2380GAT(757) ,
  \6216GAT(2411)  = ~\6207GAT(2404)  & ~\6211GAT(2407) ,
  \5507GAT(2094)  = ~\5451GAT(2068)  & ~\5450GAT(2067) ,
  \5070GAT(1927)  = ~\4891GAT(1849)  & ~\5013GAT(1900) ,
  \5613GAT(2163)  = ~\5544GAT(2134)  & ~\5370GAT(2057) ,
  \2477GAT(823)  = ~\555GAT(283)  & ~\2414GAT(782) ,
  \3715GAT(1338)  = ~\3669GAT(1319)  & ~\3668GAT(1309) ,
  \3985GAT(1434)  = ~\1050GAT(118)  & ~\3926GAT(1420) ,
  \4077GAT(1482)  = ~\4022GAT(1464)  & ~\3977GAT(1431) ,
  \2838GAT(948)  = ~\2769GAT(919)  & ~\2619GAT(852) ,
  \5404GAT(2052)  = ~\1065GAT(113)  & ~\5345GAT(2016) ,
  \723GAT(227)  = \477GAT(28)  & \52GAT(3) ,
  \1723GAT(481)  = ~\1691GAT(464)  & ~\1690GAT(463) ,
  \1693GAT(462)  = ~\1523GAT(396)  & ~\1640GAT(436) ,
  \4889GAT(1840)  = ~\4825GAT(1819)  & ~\4766GAT(1792) ,
  \1771GAT(498)  = ~\645GAT(253)  & ~\1723GAT(481) ,
  \6106GAT(2361)  = ~\6085GAT(2355)  & ~\6061GAT(2344) ,
  \4364GAT(1617)  = ~\4200GAT(1540)  & ~\4314GAT(1589) ,
  \5516GAT(2092)  = ~\5455GAT(2079)  & ~\5283GAT(1985) ,
  \6175GAT(2390)  = ~\6171GAT(2387)  & ~\6120GAT(2356) ,
  \1494GAT(350)  = ~\1122GAT(94)  & ~\1437GAT(335) ,
  \6145GAT(2375)  = ~\6141GAT(2373)  & ~\6138GAT(2372) ,
  \5621GAT(2153)  = ~\5553GAT(2132)  & ~\5552GAT(2127) ,
  \2561GAT(835)  = ~\2502GAT(811)  & ~\2501GAT(801) ,
  \1367GAT(288)  = ~\1263GAT(47) ,
  \5658GAT(2141)  = ~\5590GAT(2129)  & ~\5528GAT(2087) ,
  \1891GAT(504)  = ~\1815GAT(487)  & ~\1680GAT(426) ,
  \645GAT(253)  = \307GAT(18)  & \35GAT(2) ,
  \891GAT(171)  = \341GAT(20)  & \120GAT(7) ,
  \4943GAT(1822)  = ~\4875GAT(1813)  & ~\4704GAT(1725) ,
  \3998GAT(1424)  = ~\3943GAT(1405)  & ~\3942GAT(1404) ,
  \3043GAT(1044)  = ~\2998GAT(1025)  & ~\2997GAT(1016) ,
  \1416GAT(342)  = ~\1382GAT(321)  & ~\1381GAT(322) ,
  \4486GAT(1659)  = ~\4423GAT(1645)  & ~\4365GAT(1606) ,
  \1955GAT(575)  = ~\1836GAT(537)  & ~\1908GAT(558) ,
  \1692GAT(461)  = ~\1640GAT(436)  & ~\1591GAT(419) ,
  \5082GAT(1915)  = ~\5026GAT(1897)  & ~\4845GAT(1809) ,
  \1890GAT(506)  = ~\1173GAT(77)  & ~\1815GAT(487) ,
  \1372GAT(331)  = ~\1311GAT(302) ,
  \927GAT(159)  = \273GAT(16)  & \137GAT(8) ,
  \5235GAT(1969)  = ~\1257GAT(49)  & ~\5172GAT(1945) ,
  \3028GAT(1050)  = ~\2988GAT(1031)  & ~\2987GAT(1026) ,
  \6001GAT(2299)  = ~\5913GAT(2263)  & ~\5962GAT(2280) ,
  \6129GAT(2366)  = ~\6091GAT(2352)  & ~\6114GAT(2359) ,
  \1841GAT(534)  = ~\1775GAT(497)  & ~\1640GAT(436) ,
  \5946GAT(2286)  = ~\5846GAT(2250)  & ~\5898GAT(2268) ,
  \1854GAT(523)  = ~\1787GAT(494)  & ~\1735GAT(477) ,
  \2836GAT(937)  = ~\2769GAT(919)  & ~\2712GAT(900) ,
  \4179GAT(1549)  = ~\618GAT(262)  & ~\4114GAT(1515) ,
  \4265GAT(1561)  = ~\4140GAT(1505)  & ~\4211GAT(1527) ,
  \4098GAT(1475)  = ~\4043GAT(1457)  & ~\3998GAT(1424) ,
  \786GAT(206)  = \290GAT(17)  & \86GAT(5) ,
  \2019GAT(592)  = ~\1861GAT(522)  & ~\1975GAT(570) ,
  \2211GAT(647)  = ~\2133GAT(628)  & ~\1995GAT(565) ,
  \1032GAT(124)  = \324GAT(19)  & \171GAT(10) ,
  \4894GAT(1838)  = ~\4829GAT(1818)  & ~\4769GAT(1791) ,
  \5934GAT(2294)  = ~\633GAT(257)  & ~\5886GAT(2275) ,
  \735GAT(223)  = \273GAT(16)  & \69GAT(4) ,
  \4654GAT(1745)  = ~\4536GAT(1696)  & ~\4598GAT(1719) ,
  \3868GAT(1375)  = ~\3794GAT(1353)  & ~\3797GAT(1352) ,
  \3590GAT(1260)  = ~\3536GAT(1230)  & ~\3467GAT(1198) ,
  \4692GAT(1739)  = ~\1155GAT(83)  & ~\4634GAT(1704) ,
  \1905GAT(559)  = ~\1835GAT(539)  & ~\1834GAT(535) ,
  \2362GAT(763)  = ~\2327GAT(745)  & ~\2326GAT(742) ,
  \6195GAT(2400)  = ~\6191GAT(2397)  & ~\6082GAT(2337) ,
  \2769GAT(919)  = ~\846GAT(186)  & ~\2712GAT(900) ,
  \1983GAT(568)  = ~\1871GAT(516)  & ~\1929GAT(551) ,
  \4449GAT(1639)  = ~\1152GAT(84)  & ~\4389GAT(1611) ,
  \2743GAT(888)  = ~\2690GAT(859)  & ~\1278GAT(42) ,
  \2896GAT(976)  = ~\2842GAT(947)  & ~\2841GAT(935) ,
  \3709GAT(1341)  = ~\3665GAT(1321)  & ~\3664GAT(1313) ,
  \2971GAT(991)  = ~\1137GAT(89)  & ~\2914GAT(967) ,
  \4310GAT(1590)  = ~\4195GAT(1542)  & ~\4254GAT(1565) ,
  \2133GAT(628)  = ~\1128GAT(92)  & ~\2073GAT(608) ,
  \3624GAT(1290)  = ~\3506GAT(1243)  & ~\3568GAT(1267) ,
  \3935GAT(1407)  = ~\3882GAT(1380)  & ~\3881GAT(1371) ,
  \1373GAT(330)  = ~\1315GAT(301)  & ~\639GAT(255) ,
  \4198GAT(1530)  = ~\4130GAT(1511)  & ~\4067GAT(1484) ,
  \6277GAT(2439)  = ~\6271GAT(2437)  & ~\5666GAT(2138) ,
  \3409GAT(1179)  = ~\3311GAT(1133)  & ~\3356GAT(1152) ,
  \2993GAT(1020)  = ~\2938GAT(999)  & ~\2887GAT(979) ,
  \954GAT(150)  = \426GAT(25)  & \137GAT(8) ,
  \5168GAT(1932)  = ~\5053GAT(1883)  & ~\5109GAT(1906) ,
  \3119GAT(1057)  = ~\3058GAT(1045)  & ~\3007GAT(1009) ,
  \1556GAT(376)  = ~\1486GAT(352)  & ~\1431GAT(337) ,
  \2884GAT(980)  = ~\2822GAT(958)  & ~\2821GAT(946) ,
  \1938GAT(548)  = ~\1890GAT(506)  & ~\1889GAT(503) ,
  \1897GAT(501)  = ~\1821GAT(484)  & ~\1269GAT(45) ,
  \5026GAT(1897)  = ~\867GAT(179)  & ~\4965GAT(1866) ,
  \2210GAT(649)  = ~\1128GAT(92)  & ~\2133GAT(628) ,
  \3421GAT(1215)  = ~\612GAT(264)  & ~\3368GAT(1194) ,
  \5672GAT(2187)  = \[13] ,
  \4085GAT(1479)  = ~\4028GAT(1451)  & ~\4031GAT(1450) ,
  \5038GAT(1888)  = ~\4974GAT(1864)  & ~\4977GAT(1863) ,
  \1680GAT(426)  = ~\1573GAT(366)  & ~\1621GAT(409) ,
  \6280GAT(2443)  = \[29] ,
  \3176GAT(1092)  = ~\897GAT(169)  & ~\3107GAT(1062) ,
  \2930GAT(1001)  = ~\2813GAT(961)  & ~\2881GAT(981) ,
  \5959GAT(2281)  = ~\5912GAT(2272)  & ~\5911GAT(2264) ,
  \5975GAT(2307)  = ~\5935GAT(2293)  & ~\5938GAT(2288) ,
  \2430GAT(778)  = ~\747GAT(219)  & ~\2374GAT(759) ,
  \654GAT(250)  = \358GAT(21)  & \35GAT(2) ,
  \5440GAT(2071)  = ~\5383GAT(2054)  & ~\5200GAT(1965) ,
  \5400GAT(2044)  = ~\5277GAT(1987)  & ~\5339GAT(2019) ,
  \3433GAT(1212)  = ~\756GAT(216)  & ~\3377GAT(1189) ,
  \1856GAT(525)  = ~\1787GAT(494)  & ~\1652GAT(433) ,
  \576GAT(276)  = \460GAT(27)  & \1GAT(0) ,
  \3339GAT(1157)  = ~\3296GAT(1140)  & ~\3236GAT(1117) ,
  \4570GAT(1675)  = ~\4503GAT(1661)  & ~\4441GAT(1629) ,
  \1557GAT(377)  = ~\1026GAT(126)  & ~\1486GAT(352) ,
  \3520GAT(1236)  = ~\948GAT(152)  & ~\3449GAT(1208) ,
  \2545GAT(783)  = ~\2475GAT(765)  & ~\2474GAT(764) ,
  \4386GAT(1599)  = ~\4340GAT(1577)  & ~\4339GAT(1576) ,
  \1606GAT(414)  = ~\1552GAT(380)  & ~\1551GAT(379) ,
  \5651GAT(2142)  = ~\5586GAT(2116)  & ~\5585GAT(2115) ,
  \5450GAT(2067)  = ~\5395GAT(2045)  & ~\5336GAT(2020) ,
  \4934GAT(1824)  = ~\4871GAT(1801)  & ~\4870GAT(1800) ,
  \3332GAT(1172)  = ~\3162GAT(1099)  & ~\3280GAT(1144) ,
  \3288GAT(1142)  = ~\3172GAT(1093)  & ~\3230GAT(1120) ,
  \4348GAT(1574)  = ~\4290GAT(1564)  & ~\4238GAT(1517) ,
  \1513GAT(402)  = ~\1450GAT(361)  & ~\1315GAT(301) ,
  \5322GAT(2024)  = ~\5262GAT(1992)  & ~\5197GAT(1966) ,
  \3677GAT(1314)  = ~\3516GAT(1237)  & ~\3632GAT(1288) ,
  \3545GAT(1218)  = ~\3475GAT(1205)  & ~\3474GAT(1197) ,
  \1687GAT(468)  = ~\1508GAT(405)  & ~\1628GAT(439) ,
  \3669GAT(1319)  = ~\3496GAT(1247)  & ~\3616GAT(1292) ,
  \5540GAT(2135)  = ~\582GAT(274)  & ~\5480GAT(2105) ,
  \2093GAT(638)  = ~\648GAT(252)  & ~\2043GAT(620) ,
  \648GAT(252)  = \324GAT(19)  & \35GAT(2) ,
  \3245GAT(1113)  = ~\3198GAT(1074)  & ~\3197GAT(1073) ,
  \5706GAT(2174)  = ~\5650GAT(2144)  & ~\5649GAT(2143) ,
  \3736GAT(1330)  = ~\3681GAT(1312)  & ~\3527GAT(1224) ,
  \1720GAT(482)  = ~\1689GAT(466)  & ~\1688GAT(465) ,
  \2319GAT(701)  = ~\2265GAT(686)  & ~\2264GAT(685) ,
  \2160GAT(679)  = ~\648GAT(252)  & ~\2093GAT(638) ,
  \5360GAT(2012)  = ~\5298GAT(1980)  & ~\5301GAT(1979) ,
  \4972GAT(1865)  = ~\4916GAT(1844)  & ~\4851GAT(1806) ,
  \4460GAT(1623)  = ~\4401GAT(1595)  & ~\1296GAT(36) ,
  \4373GAT(1615)  = ~\957GAT(149)  & ~\4323GAT(1587) ,
  \3532GAT(1223)  = ~\3398GAT(1182)  & ~\3461GAT(1201) ,
  \4582GAT(1670)  = ~\4515GAT(1649)  & ~\4453GAT(1626) ,
  \3449GAT(1208)  = ~\948GAT(152)  & ~\3389GAT(1184) ,
  \3760GAT(1365)  = ~\567GAT(279)  & ~\3706GAT(1343) ,
  \6138GAT(2372)  = ~\6134GAT(2371)  & ~\6133GAT(2370) ,
  \3350GAT(1154)  = ~\3305GAT(1138)  & ~\3127GAT(1054) ,
  \4226GAT(1522)  = ~\4155GAT(1508)  & ~\3992GAT(1427) ,
  \4881GAT(1853)  = ~\4817GAT(1821)  & ~\4646GAT(1747) ,
  \4891GAT(1849)  = ~\4825GAT(1819)  & ~\4654GAT(1745) ,
  \2832GAT(953)  = ~\798GAT(202)  & ~\2765GAT(920) ,
  \4616GAT(1724)  = ~\960GAT(148)  & ~\4563GAT(1676) ,
  \1062GAT(114)  = \494GAT(29)  & \171GAT(10) ,
  \2544GAT(785)  = ~\2404GAT(748)  & ~\2470GAT(766) ,
  \1302GAT(34)  = \494GAT(29)  & \256GAT(15) ,
  \5624GAT(2152)  = ~\5554GAT(2126)  & ~\5557GAT(2125) ,
  \837GAT(189)  = \307GAT(18)  & \103GAT(6) ,
  \3806GAT(1348)  = ~\3747GAT(1327)  & ~\3746GAT(1326) ,
  \2454GAT(772)  = ~\1035GAT(123)  & ~\2392GAT(751) ,
  \1861GAT(522)  = ~\1791GAT(493)  & ~\1656GAT(432) ,
  \1512GAT(404)  = ~\594GAT(270)  & ~\1450GAT(361) ,
  \6201GAT(2402)  = ~\6197GAT(2399)  & ~\6058GAT(2325) ,
  \3922GAT(1412)  = ~\3794GAT(1353)  & ~\3868GAT(1375) ,
  \1995GAT(565)  = ~\1886GAT(507)  & ~\1938GAT(548) ,
  \4980GAT(1862)  = ~\4922GAT(1829)  & ~\4925GAT(1828) ,
  \4726GAT(1769)  = ~\912GAT(164)  & ~\4671GAT(1741) ,
  \1371GAT(332)  = ~\1311GAT(302)  & ~\591GAT(271) ,
  \3861GAT(1388)  = ~\903GAT(167)  & ~\3788GAT(1358) ,
  \2014GAT(593)  = ~\1967GAT(572)  & ~\1917GAT(555) ,
  \1422GAT(340)  = ~\1386GAT(317)  & ~\1385GAT(318) ,
  \1686GAT(467)  = ~\1628GAT(439)  & ~\1582GAT(422) ,
  \3586GAT(1270)  = ~\1095GAT(103)  & ~\3533GAT(1221) ,
  \1308GAT(32)  = \528GAT(31)  & \256GAT(15) ,
  \5421GAT(2037)  = ~\5298GAT(1980)  & ~\5360GAT(2012) ,
  \4260GAT(1562)  = ~\4205GAT(1538)  & ~\4208GAT(1528) ,
  \2833GAT(951)  = ~\2765GAT(920)  & ~\2615GAT(853) ,
  \3311GAT(1133)  = ~\3248GAT(1121)  & ~\3070GAT(1035) ,
  \3252GAT(1112)  = ~\3202GAT(1080)  & ~\3133GAT(1051) ,
  \3574GAT(1265)  = ~\3520GAT(1236)  & ~\3519GAT(1226) ,
  \1717GAT(483)  = ~\1687GAT(468)  & ~\1686GAT(467) ,
  \6058GAT(2325)  = ~\6031GAT(2314)  & ~\6030GAT(2313) ,
  \4184GAT(1547)  = ~\666GAT(246)  & ~\4118GAT(1514) ,
  \1908GAT(558)  = ~\1840GAT(536)  & ~\1839GAT(532) ,
  \2015GAT(596)  = ~\1851GAT(528)  & ~\1967GAT(572) ,
  \1713GAT(442)  = ~\1573GAT(366)  & ~\1680GAT(426) ,
  \2058GAT(615)  = ~\2019GAT(592)  & ~\2018GAT(589) ,
  \5616GAT(2154)  = ~\5548GAT(2133)  & ~\5486GAT(2101) ,
  \1305GAT(33)  = \511GAT(30)  & \256GAT(15) ,
  \5535GAT(2086)  = ~\5476GAT(2075)  & ~\5422GAT(2035) ,
  \1656GAT(432)  = ~\1543GAT(384)  & ~\1603GAT(415) ,
  \3751GAT(1335)  = ~\1194GAT(70)  & ~\3699GAT(1296) ,
  \1959GAT(574)  = ~\1841GAT(534)  & ~\1911GAT(557) ,
  \2697GAT(905)  = ~\2656GAT(886)  & ~\2655GAT(881) ,
  \2037GAT(622)  = ~\2005GAT(605)  & ~\2004GAT(603) ,
  \2161GAT(677)  = ~\2093GAT(638)  & ~\1955GAT(575) ,
  \4356GAT(1621)  = ~\4180GAT(1548)  & ~\4298GAT(1593) ,
  \987GAT(139)  = \341GAT(20)  & \154GAT(9) ,
  \4521GAT(1646)  = ~\4461GAT(1624)  & ~\4460GAT(1623) ,
  \4022GAT(1464)  = ~\954GAT(150)  & ~\3977GAT(1431) ,
  \1860GAT(524)  = ~\885GAT(173)  & ~\1791GAT(493) ,
  \5429GAT(2074)  = ~\5374GAT(2056)  & ~\5315GAT(2027) ,
  \4171GAT(1494)  = ~\4106GAT(1472)  & ~\1293GAT(37) ,
  \4478GAT(1664)  = ~\765GAT(213)  & ~\4417GAT(1637) ,
  \4466GAT(1667)  = ~\621GAT(261)  & ~\4408GAT(1642) ,
  \4408GAT(1642)  = ~\4356GAT(1621)  & ~\4355GAT(1613) ,
  \2318GAT(704)  = ~\2211GAT(647)  & ~\2260GAT(687) ,
  \5023GAT(1892)  = ~\4964GAT(1868)  & ~\4963GAT(1867) ,
  \1935GAT(549)  = ~\1885GAT(509)  & ~\1884GAT(505) ,
  \2690GAT(859)  = ~\2650GAT(841)  & ~\1278GAT(42) ,
  \2765GAT(920)  = ~\798GAT(202)  & ~\2709GAT(901) ,
  \5830GAT(2217)  = ~\5715GAT(2172)  & ~\5776GAT(2195) ,
  \4100GAT(1474)  = ~\4043GAT(1457)  & ~\3889GAT(1368) ,
  \1526GAT(394)  = ~\1462GAT(358)  & ~\1413GAT(343) ,
  \4850GAT(1808)  = ~\4727GAT(1759)  & ~\4787GAT(1786) ,
  \1511GAT(403)  = ~\1450GAT(361)  & ~\1404GAT(346) ,
  \1482GAT(353)  = ~\978GAT(142)  & ~\1428GAT(338) ,
  \2998GAT(1025)  = ~\2833GAT(951)  & ~\2946GAT(997) ,
  \1712GAT(441)  = ~\1680GAT(426)  & ~\1621GAT(409) ,
  \1803GAT(490)  = ~\1029GAT(125)  & ~\1747GAT(473) ,
  \4539GAT(1684)  = ~\4474GAT(1665)  & ~\4414GAT(1638) ,
  \852GAT(184)  = \392GAT(23)  & \103GAT(6) ,
  \4242GAT(1570)  = ~\4179GAT(1549)  & ~\4178GAT(1536) ,
  \1849GAT(526)  = ~\1783GAT(495)  & ~\1732GAT(478) ,
  \4193GAT(1531)  = ~\4126GAT(1512)  & ~\4064GAT(1486) ,
  \3647GAT(1281)  = ~\3586GAT(1270)  & ~\3404GAT(1180) ,
  \5163GAT(1933)  = ~\5103GAT(1908)  & ~\5106GAT(1907) ,
  \2446GAT(774)  = ~\939GAT(155)  & ~\2386GAT(755) ,
  \1689GAT(466)  = ~\1513GAT(402)  & ~\1632GAT(438) ,
  \3396GAT(1183)  = ~\3344GAT(1163)  & ~\3302GAT(1135) ,
  \3553GAT(1274)  = ~\3485GAT(1252)  & ~\3484GAT(1238) ,
  \5725GAT(2168)  = ~\5666GAT(2138)  & ~\5599GAT(2111) ,
  \4628GAT(1707)  = ~\4572GAT(1674)  & ~\4575GAT(1673) ,
  \4557GAT(1679)  = ~\4488GAT(1658)  & ~\4491GAT(1657) ,
  \5121GAT(1947)  = ~\5068GAT(1928)  & ~\5067GAT(1920) ,
  \1894GAT(502)  = ~\1820GAT(486)  & ~\1819GAT(485) ,
  \3678GAT(1303)  = ~\3637GAT(1287)  & ~\3636GAT(1284) ,
  \1932GAT(550)  = ~\1880GAT(512)  & ~\1879GAT(508) ,
  \2623GAT(851)  = ~\2513GAT(803)  & ~\2570GAT(832) ,
  \3895GAT(1423)  = \[8] ,
  \3187GAT(1084)  = ~\3115GAT(1060)  & ~\2962GAT(993) ,
  \3698GAT(1298)  = ~\3592GAT(1259)  & ~\3653GAT(1279) ,
  \3470GAT(1206)  = ~\1191GAT(71)  & ~\3410GAT(1177) ,
  \5569GAT(2131)  = ~\921GAT(161)  & ~\5507GAT(2094) ,
  \6036GAT(2336)  = ~\5930GAT(2295)  & ~\6005GAT(2324) ,
  \6210GAT(2408)  = \[22] ,
  \2843GAT(945)  = ~\2773GAT(918)  & ~\2623GAT(851) ,
  \4993GAT(1858)  = ~\4937GAT(1839)  & ~\4872GAT(1799) ,
  \2293GAT(710)  = ~\2181GAT(665)  & ~\2242GAT(693) ,
  \5215GAT(1960)  = ~\5151GAT(1950)  & ~\4980GAT(1862) ,
  \5200GAT(1965)  = ~\5136GAT(1942)  & ~\5139GAT(1941) ,
  \5130GAT(1952)  = ~\771GAT(211)  & ~\5073GAT(1917) ,
  \2016GAT(591)  = ~\1971GAT(571)  & ~\1920GAT(554) ,
  \3504GAT(1231)  = ~\3437GAT(1211)  & ~\3380GAT(1188) ,
  \1527GAT(395)  = ~\738GAT(222)  & ~\1462GAT(358) ,
  \4238GAT(1517)  = ~\4172GAT(1495)  & ~\4171GAT(1494) ,
  \4499GAT(1655)  = ~\4374GAT(1604)  & ~\4435GAT(1632) ,
  \5748GAT(2210)  = ~\825GAT(193)  & ~\5688GAT(2191) ,
  \2842GAT(947)  = ~\894GAT(170)  & ~\2773GAT(918) ,
  \6285GAT(2445)  = ~\6281GAT(2442)  & ~\5727GAT(2167) ,
  \3377GAT(1189)  = ~\3332GAT(1172)  & ~\3331GAT(1162) ,
  \5819GAT(2220)  = ~\5764GAT(2209)  & ~\5581GAT(2117) ,
  \4429GAT(1634)  = ~\4368GAT(1616)  & ~\4211GAT(1527) ,
  \4417GAT(1637)  = ~\4362GAT(1618)  & ~\4361GAT(1608) ,
  \3479GAT(1241)  = ~\3417GAT(1216)  & ~\3365GAT(1195) ,
  \5031GAT(1896)  = ~\915GAT(163)  & ~\4968GAT(1878) ,
  \5392GAT(2046)  = ~\5332GAT(2033)  & ~\5331GAT(2022) ,
  \3721GAT(1336)  = ~\3673GAT(1317)  & ~\3672GAT(1307) ,
  \4535GAT(1697)  = ~\669GAT(245)  & ~\4470GAT(1666) ,
  \5877GAT(2239)  = ~\5825GAT(2218)  & ~\5773GAT(2196) ,
  \2018GAT(589)  = ~\1975GAT(570)  & ~\1923GAT(553) ,
  \5528GAT(2087)  = ~\5472GAT(2061)  & ~\5471GAT(2060) ,
  \1711GAT(444)  = ~\1568GAT(369)  & ~\1676GAT(427) ,
  \4591GAT(1722)  = \[10] ,
  \3595GAT(1258)  = ~\3541GAT(1228)  & ~\3540GAT(1220) ,
  \5892GAT(2270)  = ~\5840GAT(2257)  & ~\5679GAT(2184) ,
  \5276GAT(2000)  = ~\966GAT(146)  & ~\5209GAT(1972) ,
  \999GAT(135)  = \409GAT(24)  & \154GAT(9) ,
  \5102GAT(1922)  = ~\1110GAT(98)  & ~\5047GAT(1895) ,
  \4146GAT(1503)  = ~\4079GAT(1481)  & ~\4082GAT(1480) ,
  \4380GAT(1602)  = ~\4329GAT(1580)  & ~\4332GAT(1579) ,
  \4269GAT(1571)  = ~\1005GAT(133)  & ~\4217GAT(1524) ,
  \1517GAT(401)  = ~\642GAT(254)  & ~\1454GAT(360) ,
  \729GAT(225)  = \511GAT(30)  & \52GAT(3) ,
  \789GAT(205)  = \307GAT(18)  & \86GAT(5) ,
  \4257GAT(1563)  = ~\4204GAT(1539)  & ~\4203GAT(1529) ,
  \4368GAT(1616)  = ~\909GAT(165)  & ~\4320GAT(1582) ,
  \5093GAT(1912)  = ~\4974GAT(1864)  & ~\5038GAT(1888) ,
  \3800GAT(1351)  = ~\3736GAT(1330)  & ~\3739GAT(1329) ,
  \5113GAT(1904)  = ~\5059GAT(1881)  & ~\4998GAT(1856) ,
  \1688GAT(465)  = ~\1632GAT(438)  & ~\1585GAT(421) ,
  \996GAT(136)  = \392GAT(23)  & \154GAT(9) ,
  \5227GAT(1955)  = ~\5168GAT(1932)  & ~\5167GAT(1931) ,
  \2739GAT(890)  = ~\2684GAT(861)  & ~\2687GAT(860) ,
  \6103GAT(2347)  = ~\6081GAT(2339)  & ~\6080GAT(2338) ,
  \2017GAT(594)  = ~\1856GAT(525)  & ~\1971GAT(571) ,
  \5694GAT(2179)  = ~\5633GAT(2160)  & ~\5446GAT(2069) ,
  \2694GAT(906)  = ~\2654GAT(887)  & ~\2653GAT(883) ,
  \6091GAT(2352)  = ~\6064GAT(2346)  & ~\5975GAT(2307) ,
  \2156GAT(680)  = ~\2089GAT(639)  & ~\1951GAT(576) ,
  \5301GAT(1979)  = ~\5235GAT(1969)  & ~\5234GAT(1954) ,
  \5852GAT(2248)  = ~\5798GAT(2227)  & ~\5801GAT(2226) ,
  \3031GAT(1049)  = ~\2990GAT(1030)  & ~\2989GAT(1024) ,
  \6230GAT(2418)  = \[24] ,
  \699GAT(235)  = \341GAT(20)  & \52GAT(3) ,
  \4687GAT(1730)  = ~\4628GAT(1707)  & ~\4575GAT(1673) ,
  \4094GAT(1487)  = ~\1149GAT(85)  & ~\4040GAT(1446) ,
  \1521GAT(397)  = ~\1458GAT(359)  & ~\1410GAT(344) ,
  \3616GAT(1292)  = ~\3496GAT(1247)  & ~\3562GAT(1271) ,
  \984GAT(140)  = \324GAT(19)  & \154GAT(9) ,
  \5718GAT(2171)  = ~\5659GAT(2157)  & ~\5658GAT(2141) ,
  \4006GAT(1471)  = ~\3827GAT(1401)  & ~\3947GAT(1443) ,
  \1038GAT(122)  = \358GAT(21)  & \171GAT(10) ,
  \2010GAT(597)  = ~\1959GAT(574)  & ~\1911GAT(557) ,
  \1710GAT(443)  = ~\1676GAT(427)  & ~\1618GAT(410) ,
  \2458GAT(771)  = ~\1083GAT(107)  & ~\2395GAT(750) ,
  \2371GAT(760)  = ~\2333GAT(741)  & ~\2332GAT(736) ,
  \1537GAT(389)  = ~\834GAT(190)  & ~\1470GAT(356) ,
  \5209GAT(1972)  = ~\966GAT(146)  & ~\5148GAT(1937) ,
  \696GAT(236)  = \324GAT(19)  & \52GAT(3) ,
  \5659GAT(2157)  = ~\1164GAT(80)  & ~\5590GAT(2129) ,
  \1516GAT(400)  = ~\1454GAT(360)  & ~\1407GAT(345) ,
  \1454GAT(360)  = ~\642GAT(254)  & ~\1407GAT(345) ,
  \3882GAT(1380)  = ~\1146GAT(86)  & ~\3809GAT(1356) ,
  \2615GAT(853)  = ~\2503GAT(809)  & ~\2564GAT(834) ,
  \4658GAT(1744)  = ~\4541GAT(1694)  & ~\4601GAT(1717) ,
  \5333GAT(2021)  = ~\5271GAT(2001)  & ~\5088GAT(1913) ,
  \3002GAT(1021)  = ~\2843GAT(945)  & ~\2954GAT(995) ,
  \3142GAT(1107)  = ~\3079GAT(1069)  & ~\2926GAT(1002) ,
  \3314GAT(1132)  = ~\3253GAT(1119)  & ~\3252GAT(1112) ,
  \5118GAT(1948)  = ~\5066GAT(1929)  & ~\5065GAT(1921) ,
  \4872GAT(1799)  = ~\4813GAT(1778)  & ~\4812GAT(1777) ,
  \1947GAT(577)  = ~\1826GAT(543)  & ~\1902GAT(560) ,
  \6156GAT(2381)  = ~\6147GAT(2374)  & ~\6151GAT(2377) ,
  \3474GAT(1197)  = ~\3413GAT(1185)  & ~\3362GAT(1149) ,
  \2926GAT(1002)  = ~\2808GAT(963)  & ~\2878GAT(982) ,
  \2155GAT(681)  = ~\600GAT(268)  & ~\2089GAT(639) ,
  \4328GAT(1586)  = ~\1005GAT(133)  & ~\4269GAT(1571) ,
  \606GAT(266)  = \358GAT(21)  & \18GAT(1) ,
  \5134GAT(1943)  = ~\5076GAT(1925)  & ~\5023GAT(1892) ,
  \6257GAT(2429)  = ~\6251GAT(2427)  & ~\5776GAT(2195) ,
  \4027GAT(1462)  = ~\1002GAT(134)  & ~\3980GAT(1435) ,
  \1522GAT(398)  = ~\690GAT(238)  & ~\1458GAT(359) ,
  \1999GAT(563)  = ~\1941GAT(547)  & ~\1894GAT(502) ,
  \5473GAT(2059)  = ~\5421GAT(2037)  & ~\5420GAT(2036) ,
  \6206GAT(2406)  = ~\6197GAT(2399)  & ~\6201GAT(2402) ,
  \3665GAT(1321)  = ~\3486GAT(1251)  & ~\3608GAT(1294) ,
  \2154GAT(675)  = ~\2089GAT(639)  & ~\2040GAT(621) ,
  \867GAT(179)  = \477GAT(28)  & \103GAT(6) ,
  \2139GAT(625)  = ~\2076GAT(611)  & ~\1941GAT(547) ,
  \834GAT(190)  = \290GAT(17)  & \103GAT(6) ,
  \6247GAT(2424)  = ~\6241GAT(2422)  & ~\5825GAT(2218) ,
  \3475GAT(1205)  = ~\1239GAT(55)  & ~\3413GAT(1185) ,
  \1558GAT(375)  = ~\1486GAT(352)  & ~\1351GAT(292) ,
  \5585GAT(2115)  = ~\5522GAT(2090)  & ~\5464GAT(2063) ,
  \5515GAT(2106)  = ~\1017GAT(129)  & ~\5455GAT(2079) ,
  \3027GAT(1004)  = ~\2923GAT(965)  & ~\2983GAT(984) ,
  \3693GAT(1299)  = ~\3647GAT(1281)  & ~\3650GAT(1280) ,
  \3058GAT(1045)  = ~\1041GAT(121)  & ~\3007GAT(1009) ,
  \3133GAT(1051)  = ~\3075GAT(1034)  & ~\3074GAT(1033) ,
  \4019GAT(1453)  = ~\3976GAT(1436)  & ~\3975GAT(1432) ,
  \2841GAT(935)  = ~\2773GAT(918)  & ~\2715GAT(898) ,
  \5810GAT(2222)  = ~\5760GAT(2201)  & ~\5759GAT(2200) ,
  \5801GAT(2226)  = ~\5748GAT(2210)  & ~\5747GAT(2205) ,
  \1536GAT(388)  = ~\1470GAT(356)  & ~\1419GAT(341) ,
  \6260GAT(2433)  = \[27] ,
  \2138GAT(627)  = ~\1176GAT(76)  & ~\2076GAT(611) ,
  \3794GAT(1353)  = ~\3730GAT(1342)  & ~\3577GAT(1264) ,
  \2853GAT(939)  = ~\2781GAT(916)  & ~\2631GAT(849) ,
  \5743GAT(2211)  = ~\777GAT(209)  & ~\5685GAT(2181) ,
  \3846GAT(1394)  = ~\759GAT(215)  & ~\3776GAT(1361) ,
  \2055GAT(616)  = ~\2017GAT(594)  & ~\2016GAT(591) ,
  \1379GAT(324)  = ~\1327GAT(298)  & ~\783GAT(207) ,
  \2934GAT(1000)  = ~\2818GAT(959)  & ~\2884GAT(980) ,
  \1941GAT(547)  = ~\1891GAT(504)  & ~\1894GAT(502) ,
  \3690GAT(1300)  = ~\3646GAT(1285)  & ~\3645GAT(1282) ,
  \4052GAT(1491)  = ~\4006GAT(1471)  & ~\4005GAT(1463) ,
  \2899GAT(975)  = ~\2847GAT(944)  & ~\2846GAT(934) ,
  \4353GAT(1614)  = ~\4294GAT(1594)  & ~\4242GAT(1570) ,
  \4733GAT(1757)  = ~\4677GAT(1734)  & ~\4680GAT(1733) ,
  \5596GAT(2112)  = ~\5531GAT(2104)  & ~\5360GAT(2012) ,
  \3724GAT(1334)  = ~\3675GAT(1316)  & ~\3674GAT(1306) ,
  \3268GAT(1147)  = ~\3147GAT(1105)  & ~\3215GAT(1126) ,
  \3413GAT(1185)  = ~\1239GAT(55)  & ~\3362GAT(1149) ,
  \4714GAT(1763)  = ~\4658GAT(1744)  & ~\4601GAT(1717) ,
  \5042GAT(1886)  = ~\4980GAT(1862)  & ~\4925GAT(1828) ,
  \6235GAT(2420)  = ~\6231GAT(2417)  & ~\5968GAT(2277) ,
  \2852GAT(941)  = ~\990GAT(138)  & ~\2781GAT(916) ,
  \1523GAT(396)  = ~\1458GAT(359)  & ~\1323GAT(299) ,
  \5379GAT(2055)  = ~\5256GAT(2002)  & ~\5318GAT(2026) ,
  \4839GAT(1811)  = ~\4775GAT(1798)  & ~\4607GAT(1714) ,
  \3335GAT(1159)  = ~\3288GAT(1142)  & ~\3230GAT(1120) ,
  \5865GAT(2244)  = ~\5813GAT(2233)  & ~\5761GAT(2199) ,
  \4444GAT(1641)  = ~\1104GAT(100)  & ~\4386GAT(1599) ,
  \5495GAT(2099)  = ~\5434GAT(2081)  & ~\5262GAT(1992) ,
  \771GAT(211)  = \477GAT(28)  & \69GAT(4) ,
  \5527GAT(2089)  = ~\5410GAT(2040)  & ~\5467GAT(2062) ,
  \3284GAT(1143)  = ~\3167GAT(1096)  & ~\3227GAT(1122) ,
  \1846GAT(531)  = ~\1779GAT(496)  & ~\1644GAT(435) ,
  \4884GAT(1841)  = ~\4821GAT(1820)  & ~\4763GAT(1793) ,
  \4562GAT(1678)  = ~\4429GAT(1634)  & ~\4494GAT(1656) ,
  \6176GAT(2391)  = ~\6167GAT(2384)  & ~\6171GAT(2387) ,
  \5945GAT(2285)  = ~\5898GAT(2268)  & ~\5849GAT(2249) ,
  \2997GAT(1016)  = ~\2946GAT(997)  & ~\2893GAT(977) ,
  \5489GAT(2109)  = ~\726GAT(226)  & ~\5431GAT(2073) ,
  \4540GAT(1695)  = ~\717GAT(229)  & ~\4474GAT(1665) ,
  \5114GAT(1905)  = ~\4995GAT(1857)  & ~\5059GAT(1881) ,
  \1636GAT(437)  = ~\1518GAT(399)  & ~\1588GAT(420) ,
  \609GAT(265)  = \375GAT(22)  & \18GAT(1) ,
  \5781GAT(2194)  = ~\5660GAT(2140)  & ~\5721GAT(2170) ,
  \3481GAT(1253)  = ~\3417GAT(1216)  & ~\3264GAT(1148) ,
  \3491GAT(1249)  = ~\3425GAT(1214)  & ~\3272GAT(1146) ,
  \1068GAT(112)  = \528GAT(31)  & \171GAT(10) ,
  \4195GAT(1542)  = ~\4126GAT(1512)  & ~\3963GAT(1439) ,
  \4701GAT(1726)  = ~\4642GAT(1716)  & ~\4641GAT(1703) ,
  \5700GAT(2177)  = ~\5639GAT(2147)  & ~\5642GAT(2146) ,
  \1378GAT(325)  = ~\1323GAT(299) ,
  \2012GAT(595)  = ~\1963GAT(573)  & ~\1914GAT(556) ,
  \1844GAT(529)  = ~\1779GAT(496)  & ~\1729GAT(479) ,
  \2297GAT(709)  = ~\2186GAT(662)  & ~\2245GAT(692) ,
  \5094GAT(1910)  = ~\5043GAT(1887)  & ~\5042GAT(1886) ,
  \2407GAT(747)  = ~\2358GAT(721)  & ~\2357GAT(718) ,
  \3445GAT(1209)  = ~\900GAT(168)  & ~\3386GAT(1186) ,
  \2683GAT(866)  = ~\1182GAT(74)  & ~\2644GAT(846) ,
  \6161GAT(2382)  = ~\6157GAT(2379)  & ~\6130GAT(2364) ,
  \1458GAT(359)  = ~\690GAT(238)  & ~\1410GAT(344) ,
  \4503GAT(1661)  = ~\1056GAT(116)  & ~\4441GAT(1629) ,
  \921GAT(161)  = \511GAT(30)  & \120GAT(7) ,
  \4759GAT(1749)  = ~\4643GAT(1702)  & ~\4704GAT(1725) ,
  \4890GAT(1850)  = ~\672GAT(244)  & ~\4825GAT(1819) ,
  \1035GAT(123)  = \341GAT(20)  & \171GAT(10) ,
  \579GAT(275)  = \477GAT(28)  & \1GAT(0) ,
  \2013GAT(598)  = ~\1846GAT(531)  & ~\1963GAT(573) ,
  \2567GAT(833)  = ~\2512GAT(805)  & ~\2511GAT(795) ,
  \6146GAT(2376)  = ~\6141GAT(2373) ,
  \5786GAT(2237)  = ~\5608GAT(2165)  & ~\5730GAT(2214) ,
  \5364GAT(2010)  = ~\5304GAT(1978)  & ~\1305GAT(33) ,
  \6134GAT(2371)  = ~\6108GAT(2362)  & ~\6124GAT(2367) ,
  \2205GAT(652)  = ~\1080GAT(108)  & ~\2129GAT(629) ,
  \5857GAT(2247)  = ~\5749GAT(2204)  & ~\5804GAT(2225) ,
  \1498GAT(349)  = ~\1170GAT(78)  & ~\1440GAT(334) ,
  \5988GAT(2303)  = ~\5950GAT(2292)  & ~\5904GAT(2265) ,
  \5146GAT(1938)  = ~\5088GAT(1913)  & ~\5035GAT(1889) ,
  \5663GAT(2139)  = ~\5595GAT(2128)  & ~\5594GAT(2113) ,
  \4911GAT(1832)  = ~\4845GAT(1809)  & ~\4784GAT(1787) ,
  \6009GAT(2320)  = ~\5975GAT(2307)  & ~\5938GAT(2288) ,
  \2322GAT(703)  = ~\1227GAT(59)  & ~\2266GAT(684) ,
  \864GAT(180)  = \460GAT(27)  & \103GAT(6) ,
  \6094GAT(2351)  = ~\6069GAT(2345)  & ~\6068GAT(2343) ,
  \5773GAT(2196)  = ~\5714GAT(2188)  & ~\5713GAT(2173) ,
  \4584GAT(1669)  = ~\4520GAT(1648)  & ~\4519GAT(1647) ,
  \3208GAT(1070)  = ~\3136GAT(1058)  & ~\2983GAT(984) ,
  \3657GAT(1277)  = ~\3598GAT(1257)  & ~\3545GAT(1218) ,
  \6044GAT(2331)  = ~\6014GAT(2322)  & ~\5981GAT(2304) ,
  \4808GAT(1779)  = ~\4748GAT(1752)  & ~\4751GAT(1751) ,
  \2206GAT(650)  = ~\2129GAT(629)  & ~\1991GAT(566) ,
  \4188GAT(1532)  = ~\4122GAT(1513)  & ~\4061GAT(1488) ,
  \4667GAT(1742)  = ~\4551GAT(1690)  & ~\4607GAT(1714) ,
  \2564GAT(834)  = ~\2507GAT(808)  & ~\2506GAT(798) ,
  \3938GAT(1406)  = ~\3883GAT(1370)  & ~\3886GAT(1369) ,
  \4763GAT(1793)  = ~\4711GAT(1774)  & ~\4710GAT(1766) ,
  \4010GAT(1469)  = ~\3837GAT(1397)  & ~\3955GAT(1441) ,
  \3742GAT(1328)  = ~\3687GAT(1301)  & ~\3690GAT(1300) ,
  \2773GAT(918)  = ~\894GAT(170)  & ~\2715GAT(898) ,
  \5962GAT(2280)  = ~\5913GAT(2263)  & ~\5916GAT(2262) ,
  \5256GAT(2002)  = ~\5188GAT(1974)  & ~\5017GAT(1899) ,
  \4323GAT(1587)  = ~\957GAT(149)  & ~\4266GAT(1559) ,
  \3641GAT(1286)  = ~\1047GAT(119)  & ~\3583GAT(1261) ,
  \4274GAT(1569)  = ~\1053GAT(117)  & ~\4220GAT(1535) ,
  \3152GAT(1103)  = ~\3087GAT(1067)  & ~\2934GAT(1000) ,
  \3175GAT(1081)  = ~\3107GAT(1062)  & ~\3049GAT(1041) ,
  \2851GAT(933)  = ~\2781GAT(916)  & ~\2721GAT(895) ,
  \3365GAT(1195)  = ~\3324GAT(1176)  & ~\3323GAT(1170) ,
  \6181GAT(2392)  = ~\6177GAT(2389)  & ~\6103GAT(2347) ,
  \5834GAT(2253)  = ~\5786GAT(2237)  & ~\5785GAT(2231) ,
  \4713GAT(1773)  = ~\4536GAT(1696)  & ~\4654GAT(1745) ,
  \6118GAT(2357)  = ~\6097GAT(2350)  & ~\6073GAT(2341) ,
  \4632GAT(1705)  = ~\4578GAT(1672)  & ~\4512GAT(1650) ,
  \2682GAT(862)  = ~\2644GAT(846)  & ~\2588GAT(824) ,
  \4986GAT(1859)  = ~\4933GAT(1826)  & ~\4932GAT(1825) ,
  \2619GAT(852)  = ~\2508GAT(806)  & ~\2567GAT(833) ,
  \2736GAT(891)  = ~\2683GAT(866)  & ~\2682GAT(862) ,
  \3963GAT(1439)  = ~\3847GAT(1393)  & ~\3908GAT(1416) ,
  \3171GAT(1095)  = ~\849GAT(185)  & ~\3103GAT(1063) ,
  \2217GAT(643)  = ~\2139GAT(625)  & ~\2142GAT(624) ,
  \1951GAT(576)  = ~\1831GAT(540)  & ~\1905GAT(559) ,
  \5387GAT(2048)  = ~\5327GAT(2034)  & ~\5268GAT(1989) ,
  \5443GAT(2070)  = ~\5388GAT(2053)  & ~\5387GAT(2048) ,
  \5292GAT(1998)  = ~\1161GAT(81)  & ~\5227GAT(1955) ,
  \5950GAT(2292)  = ~\828GAT(192)  & ~\5904GAT(2265) ,
  \1490GAT(351)  = ~\1074GAT(110)  & ~\1434GAT(336) ,
  \4738GAT(1756)  = ~\4622GAT(1709)  & ~\4683GAT(1732) ,
  \1591GAT(419)  = ~\1527GAT(395)  & ~\1526GAT(394) ,
  \3348GAT(1155)  = ~\3305GAT(1138)  & ~\3245GAT(1113) ,
  \4937GAT(1839)  = ~\1206GAT(66)  & ~\4872GAT(1799) ,
  \1363GAT(289)  = ~\1215GAT(63) ,
  \5431GAT(2073)  = ~\5379GAT(2055)  & ~\5378GAT(2050) ,
  \1375GAT(328)  = ~\1319GAT(300)  & ~\687GAT(239) ,
  \3971GAT(1437)  = ~\3857GAT(1389)  & ~\3914GAT(1414) ,
  \6265GAT(2435)  = ~\6261GAT(2432)  & ~\5831GAT(2215) ,
  \3383GAT(1187)  = ~\3336GAT(1169)  & ~\3335GAT(1159) ,
  \3548GAT(1217)  = ~\3476GAT(1196)  & ~\1287GAT(39) ,
  \5602GAT(2110)  = ~\5537GAT(2085)  & ~\1308GAT(32) ,
  \3292GAT(1141)  = ~\3177GAT(1090)  & ~\3233GAT(1118) ,
  \4286GAT(1554)  = ~\4161GAT(1498)  & ~\4232GAT(1520) ,
  \2552GAT(838)  = ~\2487GAT(819)  & ~\2486GAT(810) ,
  \2194GAT(651)  = ~\2121GAT(631)  & ~\2064GAT(613) ,
  \4372GAT(1605)  = ~\4323GAT(1587)  & ~\4266GAT(1559) ,
  \2121GAT(631)  = ~\984GAT(140)  & ~\2064GAT(613) ,
  \1428GAT(338)  = ~\1390GAT(313)  & ~\1389GAT(314) ,
  \2607GAT(855)  = ~\2493GAT(815)  & ~\2558GAT(836) ,
  \5565GAT(2123)  = ~\5440GAT(2071)  & ~\5501GAT(2097) ,
  \4959GAT(1869)  = ~\4901GAT(1845)  & ~\4904GAT(1835) ,
  \4721GAT(1770)  = ~\864GAT(180)  & ~\4668GAT(1736) ,
  \3674GAT(1306)  = ~\3628GAT(1289)  & ~\3571GAT(1266) ,
  \1869GAT(514)  = ~\1799GAT(491)  & ~\1744GAT(474) ,
  \2675GAT(863)  = ~\2640GAT(847)  & ~\2639GAT(844) ,
  \5578GAT(2118)  = ~\5515GAT(2106)  & ~\5514GAT(2093) ,
  \4204GAT(1539)  = ~\858GAT(182)  & ~\4134GAT(1510) ,
  \2543GAT(784)  = ~\2470GAT(766)  & ~\2407GAT(747) ,
  \2881GAT(981)  = ~\2817GAT(960)  & ~\2816GAT(949) ,
  \4047GAT(1445)  = ~\4001GAT(1433)  & ~\3944GAT(1403) ,
  \1901GAT(561)  = \[2] ,
  \1845GAT(533)  = ~\741GAT(221)  & ~\1779GAT(496) ,
  \4675GAT(1735)  = ~\4616GAT(1724)  & ~\4563GAT(1676) ,
  \4401GAT(1595)  = ~\4350GAT(1573)  & ~\1296GAT(36) ,
  \5370GAT(2057)  = ~\5246GAT(2006)  & ~\5312GAT(2028) ,
  \5768GAT(2198)  = ~\5709GAT(2189)  & ~\5651GAT(2142) ,
  \5493GAT(2100)  = ~\5434GAT(2081)  & ~\5380GAT(2049) ,
  \5088GAT(1913)  = ~\5032GAT(1890)  & ~\5035GAT(1889) ,
  \5912GAT(2272)  = ~\924GAT(160)  & ~\5861GAT(2255) ,
  \2404GAT(748)  = ~\2353GAT(723)  & ~\2217GAT(643) ,
  \567GAT(279)  = \409GAT(24)  & \1GAT(0) ,
  \726GAT(226)  = \494GAT(29)  & \52GAT(3) ,
  \3788GAT(1358)  = ~\903GAT(167)  & ~\3727GAT(1332) ,
  \4039GAT(1448)  = ~\3932GAT(1408)  & ~\3992GAT(1427) ,
  \2195GAT(658)  = ~\984GAT(140)  & ~\2121GAT(631) ,
  \5246GAT(2006)  = ~\5180GAT(1976)  & ~\5009GAT(1901) ,
  \3531GAT(1222)  = ~\3461GAT(1201)  & ~\3401GAT(1181) ,
  \1374GAT(329)  = ~\1315GAT(301) ,
  \957GAT(149)  = \443GAT(26)  & \137GAT(8) ,
  \642GAT(254)  = \290GAT(17)  & \35GAT(2) ,
  \4138GAT(1506)  = ~\4073GAT(1493)  & ~\4019GAT(1453) ,
  \831GAT(191)  = \273GAT(16)  & \103GAT(6) ,
  \6123GAT(2368)  = \[15] ,
  \5557GAT(2125)  = ~\5494GAT(2108)  & ~\5493GAT(2100) ,
  \5714GAT(2188)  = ~\1116GAT(96)  & ~\5654GAT(2158) ,
  \6111GAT(2360)  = ~\6090GAT(2354)  & ~\6089GAT(2353) ,
  \4134GAT(1510)  = ~\858GAT(182)  & ~\4070GAT(1483) ,
  \3686GAT(1310)  = ~\1047GAT(119)  & ~\3641GAT(1286) ,
  \3862GAT(1386)  = ~\3788GAT(1358)  & ~\3632GAT(1288) ,
  \3992GAT(1427)  = ~\3932GAT(1408)  & ~\3935GAT(1407) ,
  \2159GAT(672)  = ~\2093GAT(638)  & ~\2043GAT(620) ,
  \4190GAT(1544)  = ~\4122GAT(1513)  & ~\3959GAT(1440) ,
  \3856GAT(1390)  = ~\855GAT(183)  & ~\3784GAT(1359) ,
  \5629GAT(2151)  = ~\5495GAT(2099)  & ~\5560GAT(2124) ,
  \3455GAT(1203)  = ~\3392GAT(1192)  & ~\3239GAT(1116) ,
  \2386GAT(755)  = ~\2343GAT(731)  & ~\2342GAT(726) ,
  \4751GAT(1751)  = ~\4697GAT(1738)  & ~\4696GAT(1728) ,
  \3889GAT(1368)  = ~\3815GAT(1346)  & ~\3818GAT(1345) ,
  \3638GAT(1283)  = ~\3582GAT(1263)  & ~\3581GAT(1262) ,
  \5981GAT(2304)  = ~\5946GAT(2286)  & ~\5945GAT(2285) ,
  \5776GAT(2195)  = ~\5715GAT(2172)  & ~\5718GAT(2171) ,
  \2137GAT(626)  = ~\2076GAT(611)  & ~\2030GAT(578) ,
  \1685GAT(425)  = ~\1578GAT(363)  & ~\1624GAT(408) ,
  \1041GAT(121)  = \375GAT(22)  & \171GAT(10) ,
  \2403GAT(752)  = ~\1179GAT(75)  & ~\2353GAT(723) ,
  \3663GAT(1322)  = ~\3481GAT(1253)  & ~\3604GAT(1295) ,
  \3362GAT(1149)  = ~\3322GAT(1130)  & ~\3321GAT(1129) ,
  \5903GAT(2267)  = ~\5798GAT(2227)  & ~\5852GAT(2248) ,
  \5769GAT(2208)  = ~\1068GAT(112)  & ~\5709GAT(2189) ,
  \4747GAT(1765)  = ~\1155GAT(83)  & ~\4692GAT(1739) ,
  \657GAT(249)  = \375GAT(22)  & \35GAT(2) ,
  \1767GAT(499)  = ~\597GAT(269)  & ~\1720GAT(482) ,
  \5156GAT(1949)  = ~\1062GAT(114)  & ~\5097GAT(1923) ,
  \2806GAT(955)  = ~\2745GAT(925)  & ~\2694GAT(906) ,
  \6271GAT(2437)  = ~\6267GAT(2434)  & ~\5782GAT(2192) ,
  \2988GAT(1031)  = ~\2808GAT(963)  & ~\2926GAT(1002) ,
  \3840GAT(1383)  = ~\3772GAT(1362)  & ~\3715GAT(1338) ,
  \2807GAT(964)  = ~\558GAT(282)  & ~\2745GAT(925) ,
  \4103GAT(1473)  = ~\4048GAT(1455)  & ~\4047GAT(1445) ,
  \3327GAT(1166)  = ~\3272GAT(1146)  & ~\3218GAT(1125) ,
  \2196GAT(656)  = ~\2121GAT(631)  & ~\1983GAT(568) ,
  \5666GAT(2138)  = ~\5596GAT(2112)  & ~\5599GAT(2111) ,
  \1377GAT(326)  = ~\1323GAT(299)  & ~\735GAT(223) ,
  \4550GAT(1691)  = ~\813GAT(197)  & ~\4482GAT(1663) ,
  \2893GAT(977)  = ~\2837GAT(950)  & ~\2836GAT(937) ,
  \5172GAT(1945)  = ~\1257GAT(49)  & ~\5115GAT(1903) ,
  \2674GAT(870)  = ~\2528GAT(794)  & ~\2635GAT(848) ,
  \5789GAT(2229)  = ~\5739GAT(2212)  & ~\5738GAT(2207) ,
  \3730GAT(1342)  = ~\951GAT(151)  & ~\3678GAT(1303) ,
  \3207GAT(1078)  = ~\1236GAT(56)  & ~\3136GAT(1058) ,
  \4534GAT(1685)  = ~\4470GAT(1666)  & ~\4411GAT(1640) ,
  \4151GAT(1502)  = ~\4028GAT(1451)  & ~\4085GAT(1479) ,
  \4611GAT(1712)  = ~\4557GAT(1679)  & ~\4491GAT(1657) ,
  \2332GAT(736)  = ~\2281GAT(713)  & ~\2233GAT(696) ,
  \1553GAT(378)  = ~\1482GAT(353)  & ~\1347GAT(293) ,
  \5630GAT(2149)  = ~\5565GAT(2123)  & ~\5564GAT(2122) ,
  \951GAT(151)  = \409GAT(24)  & \137GAT(8) ,
  \4662GAT(1743)  = ~\4546GAT(1692)  & ~\4604GAT(1715) ,
  \1538GAT(387)  = ~\1470GAT(356)  & ~\1335GAT(296) ,
  \1967GAT(572)  = ~\1851GAT(528)  & ~\1917GAT(555) ,
  \1065GAT(113)  = \511GAT(30)  & \171GAT(10) ,
  \6227GAT(2414)  = ~\6221GAT(2412)  & ~\5919GAT(2261) ,
  \4355GAT(1613)  = ~\4298GAT(1593)  & ~\4245GAT(1568) ,
  \5067GAT(1920)  = ~\5009GAT(1901)  & ~\4950GAT(1873) ,
  \4164GAT(1497)  = ~\4099GAT(1485)  & ~\4098GAT(1475) ,
  \5590GAT(2129)  = ~\1164GAT(80)  & ~\5528GAT(2087) ,
  \2214GAT(644)  = ~\2138GAT(627)  & ~\2137GAT(626) ,
  \1747GAT(473)  = ~\1707GAT(448)  & ~\1706GAT(447) ,
  \4183GAT(1534)  = ~\4118GAT(1514)  & ~\4058GAT(1489) ,
  \3121GAT(1056)  = ~\3058GAT(1045)  & ~\2908GAT(970) ,
  \1684GAT(424)  = ~\1624GAT(408)  & ~\1266GAT(46) ,
  \3792GAT(1354)  = ~\3730GAT(1342)  & ~\3678GAT(1303) ,
  \5160GAT(1934)  = ~\5102GAT(1922)  & ~\5101GAT(1909) ,
  \2333GAT(741)  = ~\2166GAT(674)  & ~\2281GAT(713) ,
  \4625GAT(1708)  = ~\4571GAT(1687)  & ~\4570GAT(1675) ,
  \1864GAT(517)  = ~\1795GAT(492)  & ~\1741GAT(475) ,
  \3429GAT(1213)  = ~\708GAT(232)  & ~\3374GAT(1191) ,
  \3301GAT(1139)  = ~\3187GAT(1084)  & ~\3239GAT(1116) ,
  \5798GAT(2227)  = ~\5743GAT(2211)  & ~\5560GAT(2124) ,
  \1251GAT(51)  = \477GAT(28)  & \239GAT(14) ,
  \1431GAT(337)  = ~\1392GAT(311)  & ~\1391GAT(312) ,
  \1552GAT(380)  = ~\978GAT(142)  & ~\1482GAT(353) ,
  \2731GAT(893)  = ~\2678GAT(868)  & ~\2641GAT(843) ,
  \5205GAT(1964)  = ~\5082GAT(1915)  & ~\5142GAT(1940) ,
  \1376GAT(327)  = ~\1319GAT(300) ,
  \2097GAT(637)  = ~\696GAT(236)  & ~\2046GAT(619) ,
  \2890GAT(978)  = ~\2832GAT(953)  & ~\2831GAT(940) ,
  \1254GAT(50)  = \494GAT(29)  & \239GAT(14) ,
  \4001GAT(1433)  = ~\1245GAT(53)  & ~\3944GAT(1403) ,
  \4441GAT(1629)  = ~\4385GAT(1601)  & ~\4384GAT(1600) ,
  \3827GAT(1401)  = ~\3760GAT(1365)  & ~\3604GAT(1295) ,
  \1865GAT(521)  = ~\933GAT(157)  & ~\1795GAT(492) ,
  \2803GAT(907)  = ~\2744GAT(889)  & ~\2743GAT(888) ,
  \651GAT(251)  = \341GAT(20)  & \35GAT(2) ,
  \2732GAT(897)  = ~\1134GAT(90)  & ~\2678GAT(868) ,
  \1991GAT(566)  = ~\1881GAT(510)  & ~\1935GAT(549) ,
  \5135GAT(1951)  = ~\819GAT(195)  & ~\5076GAT(1925) ,
  \3182GAT(1087)  = ~\3111GAT(1061)  & ~\2958GAT(994) ,
  \2248GAT(691)  = ~\2195GAT(658)  & ~\2194GAT(651) ,
  \564GAT(280)  = \392GAT(23)  & \1GAT(0) ,
  \3276GAT(1145)  = ~\3157GAT(1101)  & ~\3221GAT(1124) ,
  \5739GAT(2212)  = ~\5618GAT(2161)  & ~\5679GAT(2184) ,
  \6215GAT(2410)  = ~\6211GAT(2407)  & ~\6032GAT(2312) ,
  \3328GAT(1174)  = ~\3152GAT(1103)  & ~\3272GAT(1146) ,
  \5244GAT(1997)  = ~\5180GAT(1976)  & ~\5121GAT(1947) ,
  \6170GAT(2388)  = \[18] ,
  \573GAT(277)  = \443GAT(26)  & \1GAT(0) ,
  \5142GAT(1940)  = ~\5082GAT(1915)  & ~\5085GAT(1914) ,
  \5891GAT(2274)  = ~\681GAT(241)  & ~\5840GAT(2257) ,
  \3598GAT(1257)  = ~\3542GAT(1219)  & ~\3545GAT(1218) ,
  \6107GAT(2363)  = ~\588GAT(272)  & ~\6085GAT(2355) ,
  \5408GAT(2041)  = ~\5348GAT(2032)  & ~\5289GAT(1982) ,
  \2450GAT(773)  = ~\987GAT(139)  & ~\2389GAT(753) ,
  \3006GAT(1017)  = ~\2853GAT(939)  & ~\2962GAT(993) ,
  \3341GAT(1156)  = ~\3301GAT(1139)  & ~\3300GAT(1136) ,
  \1744GAT(474)  = ~\1705GAT(450)  & ~\1704GAT(449) ,
  \2329GAT(744)  = ~\2156GAT(680)  & ~\2273GAT(715) ,
  \3264GAT(1148)  = ~\3142GAT(1107)  & ~\3212GAT(1127) ,
  \5761GAT(2199)  = ~\5705GAT(2176)  & ~\5704GAT(2175) ,
  \936GAT(156)  = \324GAT(19)  & \137GAT(8) ,
  \4015GAT(1456)  = ~\3967GAT(1438)  & ~\3911GAT(1415) ,
  \5271GAT(2001)  = ~\918GAT(162)  & ~\5206GAT(1962) ,
  \3976GAT(1436)  = ~\3862GAT(1386)  & ~\3917GAT(1413) ,
  \1902GAT(560)  = ~\1830GAT(542)  & ~\1829GAT(538) ,
  \777GAT(209)  = \511GAT(30)  & \69GAT(4) ,
  \5955GAT(2291)  = ~\876GAT(176)  & ~\5907GAT(2273) ,
  \3386GAT(1186)  = ~\3338GAT(1167)  & ~\3337GAT(1158) ,
  \4281GAT(1555)  = ~\4226GAT(1522)  & ~\4229GAT(1521) ,
  \3951GAT(1442)  = ~\3832GAT(1399)  & ~\3899GAT(1421) ,
  \3243GAT(1114)  = ~\3193GAT(1075)  & ~\3124GAT(1055) ,
  \2027GAT(584)  = ~\1881GAT(510)  & ~\1991GAT(566) ,
  \4637GAT(1718)  = ~\1203GAT(67)  & ~\4584GAT(1669) ,
  \4718GAT(1761)  = ~\4667GAT(1742)  & ~\4666GAT(1737) ,
  \6288GAT(2447)  = \[31] ,
  \4494GAT(1656)  = ~\4429GAT(1634)  & ~\4432GAT(1633) ,
  \3984GAT(1430)  = ~\3926GAT(1420)  & ~\3874GAT(1372) ,
  \4974GAT(1864)  = ~\4916GAT(1844)  & ~\4733GAT(1757) ,
  \4942GAT(1837)  = ~\1254GAT(50)  & ~\4875GAT(1813) ,
  \5548GAT(2133)  = ~\678GAT(242)  & ~\5486GAT(2101) ,
  \3814GAT(1355)  = ~\1194GAT(70)  & ~\3751GAT(1335) ,
  \5506GAT(2096)  = ~\5389GAT(2047)  & ~\5446GAT(2069) ,
  \4592GAT(1721)  = ~\4530GAT(1699)  & ~\4529GAT(1686) ,
  \5929GAT(2296)  = ~\585GAT(273)  & ~\5882GAT(2276) ,
  \5059GAT(1881)  = ~\4995GAT(1857)  & ~\4998GAT(1856) ,
  \3893GAT(1366)  = ~\3821GAT(1344)  & ~\1290GAT(38) ,
  \6276GAT(2441)  = ~\6267GAT(2434)  & ~\6271GAT(2437) ,
  \4254GAT(1565)  = ~\4199GAT(1541)  & ~\4198GAT(1530) ,
  \3671GAT(1318)  = ~\3501GAT(1245)  & ~\3620GAT(1291) ,
  \2802GAT(909)  = ~\2684GAT(861)  & ~\2739GAT(890) ,
  \5760GAT(2201)  = ~\5639GAT(2147)  & ~\5700GAT(2177) ,
  \3490GAT(1250)  = ~\660GAT(248)  & ~\3425GAT(1214) ,
  \3083GAT(1068)  = ~\609GAT(265)  & ~\3031GAT(1049) ,
  \5822GAT(2219)  = ~\5769GAT(2208)  & ~\5768GAT(2198) ,
  \5967GAT(2279)  = ~\5867GAT(2243)  & ~\5919GAT(2261) ,
  \3768GAT(1363)  = ~\663GAT(247)  & ~\3712GAT(1339) ,
  \5752GAT(2203)  = ~\5693GAT(2190)  & ~\5692GAT(2180) ,
  \1914GAT(556)  = ~\1850GAT(530)  & ~\1849GAT(526) ,
  \2330GAT(738)  = ~\2277GAT(714)  & ~\2230GAT(697) ,
  \2328GAT(740)  = ~\2273GAT(715)  & ~\2227GAT(698) ,
  \570GAT(278)  = \426GAT(25)  & \1GAT(0) ,
  \5309GAT(2029)  = ~\5245GAT(2007)  & ~\5244GAT(1997) ,
  \636GAT(256)  = \528GAT(31)  & \18GAT(1) ,
  \4340GAT(1577)  = ~\4226GAT(1522)  & ~\4281GAT(1555) ,
  \1551GAT(379)  = ~\1482GAT(353)  & ~\1428GAT(338) ,
  \4199GAT(1541)  = ~\810GAT(198)  & ~\4130GAT(1511) ,
  \4515GAT(1649)  = ~\4450GAT(1627)  & ~\4453GAT(1626) ,
  \5001GAT(1855)  = ~\4943GAT(1822)  & ~\1302GAT(34) ,
  \2026GAT(581)  = ~\1991GAT(566)  & ~\1935GAT(549) ,
  \2848GAT(942)  = ~\2777GAT(917)  & ~\2627GAT(850) ,
  \5574GAT(2130)  = ~\969GAT(145)  & ~\5510GAT(2107) ,
  \6000GAT(2298)  = ~\5962GAT(2280)  & ~\5916GAT(2262) ,
  \3877GAT(1382)  = ~\1098GAT(102)  & ~\3806GAT(1348) ,
  \5649GAT(2143)  = ~\5581GAT(2117)  & ~\5519GAT(2091) ,
  \3218GAT(1125)  = ~\3156GAT(1102)  & ~\3155GAT(1088) ,
  \5236GAT(1953)  = ~\5172GAT(1945)  & ~\5001GAT(1855) ,
  \801GAT(201)  = \375GAT(22)  & \86GAT(5) ,
  \5904GAT(2265)  = ~\5857GAT(2247)  & ~\5856GAT(2246) ,
  \2389GAT(753)  = ~\2345GAT(729)  & ~\2344GAT(724) ,
  \2817GAT(960)  = ~\654GAT(250)  & ~\2753GAT(923) ,
  \5071GAT(1918)  = ~\5017GAT(1899)  & ~\4956GAT(1870) ,
  \2082GAT(606)  = ~\2033GAT(580)  & ~\1897GAT(501) ,
  \3511GAT(1240)  = ~\3441GAT(1210)  & ~\3288GAT(1142) ,
  \1866GAT(519)  = ~\1795GAT(492)  & ~\1660GAT(431) ,
  \2678GAT(868)  = ~\1134GAT(90)  & ~\2641GAT(843) ,
  \5298GAT(1980)  = ~\5230GAT(1970)  & ~\5059GAT(1881) ,
  \3997GAT(1426)  = ~\3883GAT(1370)  & ~\3938GAT(1406) ,
  \6005GAT(2324)  = ~\5930GAT(2295)  & ~\5972GAT(2308) ,
  \1531GAT(391)  = ~\1466GAT(357)  & ~\1416GAT(342) ,
  \1381GAT(322)  = ~\1331GAT(297)  & ~\831GAT(191) ,
  \2129GAT(629)  = ~\1080GAT(108)  & ~\2070GAT(610) ,
  \4904GAT(1835)  = ~\4838GAT(1816)  & ~\4837GAT(1812) ,
  \2442GAT(775)  = ~\891GAT(171)  & ~\2383GAT(756) ,
  \2808GAT(963)  = ~\2745GAT(925)  & ~\2595GAT(858) ,
  \3706GAT(1343)  = ~\3663GAT(1322)  & ~\3662GAT(1315) ,
  \6080GAT(2338)  = ~\6052GAT(2328)  & ~\6023GAT(2316) ,
  \5318GAT(2026)  = ~\5256GAT(2002)  & ~\5259GAT(1993) ,
  \2733GAT(892)  = ~\2678GAT(868)  & ~\2539GAT(786) ,
  \4512GAT(1650)  = ~\4449GAT(1639)  & ~\4448GAT(1628) ,
  \963GAT(147)  = \477GAT(28)  & \137GAT(8) ,
  \711GAT(231)  = \409GAT(24)  & \52GAT(3) ,
  \2331GAT(743)  = ~\2161GAT(677)  & ~\2277GAT(714) ,
  \5103GAT(1908)  = ~\5047GAT(1895)  & ~\4866GAT(1802) ,
  \2801GAT(908)  = ~\2739GAT(890)  & ~\2687GAT(860) ,
  \2025GAT(586)  = ~\1876GAT(513)  & ~\1987GAT(567) ,
  \3776GAT(1361)  = ~\759GAT(215)  & ~\3718GAT(1337) ,
  \3344GAT(1163)  = ~\1044GAT(120)  & ~\3302GAT(1135) ,
  \5017GAT(1899)  = ~\4896GAT(1847)  & ~\4956GAT(1870) ,
  \1425GAT(339)  = ~\1388GAT(315)  & ~\1387GAT(316) ,
  \3155GAT(1088)  = ~\3091GAT(1066)  & ~\3037GAT(1047) ,
  \2846GAT(934)  = ~\2777GAT(917)  & ~\2718GAT(896) ,
  \2847GAT(944)  = ~\942GAT(154)  & ~\2777GAT(917) ,
  \6052GAT(2328)  = ~\6020GAT(2317)  & ~\6023GAT(2316) ,
  \2081GAT(609)  = ~\1224GAT(60)  & ~\2033GAT(580) ,
  \1359GAT(290)  = ~\1167GAT(79) ,
  \2327GAT(745)  = ~\2151GAT(682)  & ~\2269GAT(716) ,
  \3022GAT(1005)  = ~\2977GAT(986)  & ~\2980GAT(985) ,
  \4009GAT(1460)  = ~\3955GAT(1441)  & ~\3902GAT(1419) ,
  \4995GAT(1857)  = ~\4937GAT(1839)  & ~\4754GAT(1750) ,
  \5461GAT(2064)  = ~\5404GAT(2052)  & ~\5221GAT(1958) ,
  \2464GAT(768)  = ~\2398GAT(754)  & ~\2260GAT(687) ,
  \2858GAT(936)  = ~\2785GAT(915)  & ~\2635GAT(848) ,
  \600GAT(268)  = \324GAT(19)  & \18GAT(1) ,
  \5139GAT(1941)  = ~\5081GAT(1924)  & ~\5080GAT(1916) ,
  \1799GAT(491)  = ~\981GAT(141)  & ~\1744GAT(474) ,
  \1380GAT(323)  = ~\1327GAT(298) ,
  \4349GAT(1584)  = ~\1248GAT(52)  & ~\4290GAT(1564) ,
  \3371GAT(1193)  = ~\3328GAT(1174)  & ~\3327GAT(1166) ,
  \5692GAT(2180)  = ~\5633GAT(2160)  & ~\5566GAT(2121) ,
  \5846GAT(2250)  = ~\5792GAT(2235)  & ~\5624GAT(2152) ,
  \4742GAT(1767)  = ~\1107GAT(99)  & ~\4689GAT(1729) ,
  \5169GAT(1930)  = ~\5114GAT(1905)  & ~\5113GAT(1904) ,
  \4482GAT(1663)  = ~\813GAT(197)  & ~\4420GAT(1636) ,
  \2992GAT(1029)  = ~\2818GAT(959)  & ~\2934GAT(1000) ,
  \1566GAT(370)  = ~\1494GAT(350)  & ~\1437GAT(335) ,
  \5536GAT(2102)  = ~\1260GAT(48)  & ~\5476GAT(2075) ,
  \5673GAT(2186)  = ~\5612GAT(2164)  & ~\5611GAT(2155) ,
  \2641GAT(843)  = ~\2587GAT(826)  & ~\2586GAT(825) ,
  \2818GAT(959)  = ~\2753GAT(923)  & ~\2603GAT(856) ,
  \5068GAT(1928)  = ~\4886GAT(1851)  & ~\5009GAT(1901) ,
  \6114GAT(2359)  = ~\6091GAT(2352)  & ~\6094GAT(2351) ,
  \1071GAT(111)  = \273GAT(16)  & \188GAT(11) ,
  \4470GAT(1666)  = ~\669GAT(245)  & ~\4411GAT(1640) ,
  \4448GAT(1628)  = ~\4389GAT(1611)  & ~\4341GAT(1575) ,
  \2958GAT(994)  = ~\2848GAT(942)  & ~\2902GAT(973) ,
  \4114GAT(1515)  = ~\618GAT(262)  & ~\4055GAT(1490) ,
  \3167GAT(1096)  = ~\3099GAT(1064)  & ~\2946GAT(997) ,
  \2987GAT(1026)  = ~\2926GAT(1002)  & ~\2878GAT(982) ,
  \1532GAT(392)  = ~\786GAT(206)  & ~\1466GAT(357) ,
  \2640GAT(847)  = ~\2533GAT(791)  & ~\2582GAT(827) ,
  \4266GAT(1559)  = ~\4216GAT(1526)  & ~\4215GAT(1525) ,
  \4374GAT(1604)  = ~\4323GAT(1587)  & ~\4146GAT(1503) ,
  \3672GAT(1307)  = ~\3624GAT(1290)  & ~\3568GAT(1267) ,
  \3818GAT(1345)  = ~\3756GAT(1333)  & ~\3755GAT(1324) ,
  \5730GAT(2214)  = ~\5608GAT(2165)  & ~\5673GAT(2186) ,
  \1383GAT(320)  = ~\1335GAT(296)  & ~\879GAT(175) ,
  \5638GAT(2159)  = ~\921GAT(161)  & ~\5569GAT(2131) ,
  \3666GAT(1311)  = ~\3612GAT(1293)  & ~\3559GAT(1272) ,
  \5660GAT(2140)  = ~\5590GAT(2129)  & ~\5416GAT(2038) ,
  \4561GAT(1677)  = ~\4494GAT(1656)  & ~\4432GAT(1633) ,
  \2080GAT(607)  = ~\2033GAT(580)  & ~\2001GAT(562) ,
  \5925GAT(2258)  = ~\5878GAT(2240)  & ~\5877GAT(2239) ,
  \4796GAT(1796)  = ~\1059GAT(115)  & ~\4739GAT(1754) ;
endmodule

