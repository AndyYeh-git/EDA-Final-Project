// Benchmark "test1" written by ABC on Thu Jun 27 17:57:52 2019

module test1 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n,
    o, p, q, r, s, t, u, v  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n;
  output o, p, q, r, s, t, u, v;
  wire new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_,
    new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_,
    new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_,
    new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_;
  gate1 g000(j, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n23_);
  gate1 g001(new_n23_, i, 1'b0, 1'b0, 1'b0, 1'b1, new_n24_);
  gate1 g002(k, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n25_);
  gate1 g003(l, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n26_);
  gate1 g004(n, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n27_);
  gate1 g005(new_n27_, new_n26_, 1'b0, 1'b0, 1'b0, new_n25_, new_n28_);
  gate1 g006(n, k, 1'b0, 1'b0, 1'b0, 1'b1, new_n29_);
  gate1 g007(new_n29_, ew_n28_), .c(new_n24_, 1'b0, 1'b1, new_n28_, 1'b1, new_n30_);
  gate1 g008(a, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n31_);
  gate1 g009(e, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n32_);
  gate1 g010(new_n32_, new_n31_, 1'b0, 1'b0, 1'b0, 1'b1, new_n33_);
  gate1 g011(new_n33_, new_n30_, 1'b0, 1'b0, 1'b0, 1'b1, new_n34_);
  gate1 g012(i, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n35_);
  gate1 g013(new_n27_, new_n25_, 1'b0, 1'b0, 1'b0, new_n35_, new_n36_);
  gate1 g014(l, ), .c(new_n36_, 1'b0, 1'b1, j, 1'b1, new_n37_);
  gate1 g015(new_n37_, new_n31_, 1'b0, 1'b0, 1'b0, 1'b1, new_n38_);
  gate1 g016(n, j, 1'b0, 1'b0, 1'b0, new_n35_, new_n39_);
  gate1 g017(new_n39_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n40_);
  gate1 g018(new_n26_, k, 1'b0, 1'b0, 1'b0, 1'b1, new_n41_);
  gate1 g019(e, new_n31_, 1'b0, 1'b0, 1'b0, 1'b1, new_n42_);
  gate1 g020(new_n42_, new_n41_, 1'b0, 1'b1, 1'b1, 1'b1, new_n43_);
  gate1 g021(e, new_n31_, 1'b0, 1'b1, 1'b1, 1'b1, new_n44_);
  oai21  g022(.a(new_n44_), .b(new_n43_), .c(new_n40_), .O(new_n45_));
  gate1 g023(new_n45_, new_n38_, 1'b0, 1'b0, 1'b0, new_n34_, new_n46_);
  gate1 g024(new_n46_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n47_);
  gate1 g025(e, a, 1'b0, 1'b0, 1'b0, 1'b1, new_n48_);
  gate1 g026(new_n48_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n49_);
  gate1 g027(new_n23_, i, 1'b0, 1'b1, 1'b1, 1'b1, new_n50_);
  gate1 g028(new_n50_, new_n41_, 1'b0, 1'b0, 1'b0, n, new_n51_);
  gate1 g029(n, j, 1'b0, 1'b1, 1'b1, 1'b1, new_n52_);
  gate1 g030(k, i, 1'b1, 1'b1, 1'b1, 1'b0, new_n53_);
  gate1 g031(new_n53_, new_n52_, 1'b0, 1'b0, 1'b0, l, new_n54_);
  gate1 g032(j, i, 1'b0, 1'b0, 1'b0, 1'b1, new_n55_);
  gate1 g033(new_n55_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n56_);
  gate1 g034(new_n56_, new_n26_, 1'b0, 1'b0, 1'b0, k, new_n57_);
  gate1 g035(new_n57_, new_n54_, 1'b0, 1'b0, 1'b0, new_n51_, new_n58_);
  gate1 g036(new_n26_, k, 1'b0, 1'b0, 1'b0, new_n35_, new_n59_);
  gate1 g037(new_n59_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n60_);
  gate1 g038(new_n60_, new_n23_, 1'b0, 1'b0, 1'b0, 1'b1, new_n61_);
  gate1 g039(l, new_n25_, 1'b0, 1'b0, 1'b0, 1'b1, new_n62_);
  gate1 g040(new_n23_, new_n35_, 1'b0, 1'b0, 1'b0, 1'b1, new_n63_);
  gate1 g041(new_n63_, ew_n55_), .c(new_n62_, 1'b0, 1'b1, new_n55_, 1'b1, new_n64_);
  gate1 g042(new_n64_, n, 1'b0, 1'b0, 1'b0, 1'b1, new_n65_);
  gate1 g043(new_n65_, new_n61_, 1'b0, 1'b0, 1'b0, 1'b1, new_n66_);
  aoi22  g044(.a(new_n66_), .b(new_n49_), .c(new_n58_), .d(new_n32_), .O(new_n67_));
  gate1 g045(new_n67_, new_n47_, 1'b0, 1'b0, 1'b0, 1'b1, new_n68_);
  gate1 g046(n, j, 1'b1, 1'b1, 1'b1, 1'b0, new_n69_);
  gate1 g047(new_n69_, l, 1'b0, 1'b0, 1'b0, new_n35_, new_n70_);
  gate1 g048(new_n70_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n71_);
  gate1 g049(new_n71_, new_n49_, 1'b0, 1'b0, 1'b0, new_n25_, new_n72_);
  gate1 g050(new_n26_, k, 1'b0, 1'b0, 1'b0, i, new_n73_);
  gate1 g051(new_n73_, new_n27_, j, 1'b1, 1'b1, 1'b1, new_n74_);
  gate1 g052(n, new_n26_, 1'b0, 1'b0, 1'b0, k, new_n75_);
  gate1 g053(new_n75_, new_n55_, 1'b0, 1'b1, 1'b1, 1'b1, new_n76_);
  gate1 g054(new_n76_, new_n68_, 1'b0, 1'b0, 1'b0, a, new_n77_);
  gate1 g055(new_n58_, new_n32_, 1'b0, 1'b0, 1'b0, 1'b1, new_n78_);
  aoi22  g056(.a(new_n64_), .b(n), .c(new_n60_), .d(new_n23_), .O(new_n79_));
  oai21  g057(.a(new_n79_), .b(new_n48_), .c(new_n78_), .O(new_n80_));
  oai21  g058(.a(new_n80_), .b(new_n46_), .c(new_n71_), .O(new_n81_));
  gate1 g059(new_n75_, new_n63_, 1'b0, 1'b1, 1'b1, 1'b1, new_n82_);
  gate1 g060(new_n82_, new_n67_, 1'b0, 1'b0, 1'b0, new_n47_, new_n83_);
  gate1 g061(new_n75_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n84_);
  gate1 g062(new_n24_, new_n48_, 1'b0, 1'b1, 1'b1, 1'b1, new_n85_);
  aoi22  g063(.a(new_n85_), .b(new_n84_), .c(new_n71_), .d(a), .O(new_n86_));
  gate1 g064(new_n86_, new_n83_, 1'b0, 1'b0, 1'b0, new_n81_, new_n87_);
  gate1 g065(new_n87_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n88_);
  gate1 g066(new_n88_, new_n77_, 1'b0, 1'b0, 1'b0, new_n74_, new_n89_);
  gate1 g067(new_n89_, new_n72_, 1'b0, 1'b0, 1'b0, 1'b1, new_n90_);
  gate1 g068(new_n90_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n91_);
  gate1 g069(new_n53_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n92_);
  gate1 g070(n, new_n26_, 1'b0, 1'b0, 1'b0, new_n23_, new_n93_);
  gate1 g071(new_n93_, new_n92_, 1'b0, 1'b1, 1'b1, 1'b1, new_n94_);
  gate1 g072(new_n94_, new_n91_, 1'b0, 1'b0, 1'b0, new_n68_, new_n95_);
  gate1 g073(new_n88_, new_n77_, 1'b0, 1'b0, 1'b0, 1'b1, new_n96_);
  gate1 g074(k, new_n35_, 1'b0, 1'b0, 1'b0, new_n31_, new_n97_);
  gate1 g075(new_n97_, new_n93_, 1'b0, 1'b1, 1'b1, 1'b1, new_n98_);
  gate1 g076(new_n29_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n99_);
  gate1 g077(l, a, 1'b1, 1'b1, 1'b1, 1'b0, new_n100_);
  gate1 g078(new_n100_, new_n55_, 1'b0, 1'b0, 1'b0, new_n99_, new_n101_);
  gate1 g079(new_n101_, new_n80_, new_n46_, 1'b1, 1'b1, 1'b1, new_n102_);
  gate1 g080(new_n93_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n103_);
  gate1 g081(k, new_n35_, 1'b0, 1'b1, 1'b1, 1'b1, new_n104_);
  gate1 g082(new_n104_, new_n103_, 1'b0, 1'b0, 1'b0, e, new_n105_);
  gate1 g083(new_n32_, a, 1'b0, 1'b1, 1'b1, 1'b1, new_n106_);
  gate1 g084(new_n24_, new_n27_, k, 1'b1, 1'b1, 1'b1, new_n107_);
  oai21  g085(.a(new_n44_), .b(new_n106_), .c(new_n107_), .O(new_n108_));
  gate1 g086(k, j, 1'b0, 1'b0, 1'b0, i, new_n109_);
  gate1 g087(new_n109_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n110_);
  gate1 g088(new_n27_, new_n26_, a, 1'b1, 1'b1, 1'b1, new_n111_);
  gate1 g089(n, new_n25_, 1'b0, 1'b0, 1'b0, new_n35_, new_n112_);
  gate1 g090(new_n112_, l, new_n31_, 1'b1, 1'b1, 1'b1, new_n113_);
  gate1 g091(new_n111_, ew_n110_), .c(new_n113_, 1'b0, 1'b1, new_n110_, 1'b1, new_n114_);
  gate1 g092(new_n114_, new_n108_, 1'b0, 1'b0, 1'b0, new_n105_, new_n115_);
  gate1 g093(new_n115_, new_n102_, 1'b0, 1'b1, 1'b1, 1'b1, new_n116_);
  gate1 g094(new_n23_, a, 1'b0, 1'b0, 1'b0, 1'b1, new_n117_);
  gate1 g095(new_n117_, new_n112_, new_n68_, 1'b1, 1'b1, 1'b1, new_n118_);
  gate1 g096(new_n112_, l, new_n23_, 1'b1, 1'b1, 1'b1, new_n119_);
  gate1 g097(new_n119_, ew_n68_), .c(new_n118_, 1'b0, 1'b1, new_n68_, 1'b1, new_n120_);
  gate1 g098(n, l, 1'b0, 1'b0, 1'b0, new_n31_, new_n121_);
  gate1 g099(new_n63_, ew_n25_), .c(new_n121_, 1'b0, 1'b1, new_n25_, 1'b1, new_n122_);
  gate1 g100(new_n25_, j, 1'b0, 1'b0, 1'b0, i, new_n123_);
  oai22  g101(.a(new_n123_), .b(new_n26_), .c(new_n59_), .d(new_n23_), .O(new_n124_));
  gate1 g102(new_n124_, n, 1'b0, 1'b0, 1'b0, 1'b1, new_n125_);
  gate1 g103(new_n125_, new_n80_, new_n46_, 1'b1, 1'b1, 1'b1, new_n126_);
  gate1 g104(new_n122_, ew_n68_), .c(new_n126_, 1'b0, 1'b1, new_n68_, 1'b1, new_n127_);
  gate1 g105(new_n127_, new_n120_, 1'b0, 1'b0, 1'b0, new_n116_, new_n128_);
  gate1 g106(new_n98_, ew_n96_), .c(new_n128_, 1'b0, 1'b1, new_n96_, 1'b1, new_n129_);
  gate1 g107(new_n96_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n130_);
  gate1 g108(new_n93_, i, new_n31_, 1'b1, 1'b1, 1'b1, new_n131_);
  oai21  g109(.a(new_n131_), .b(new_n76_), .c(new_n130_), .O(new_n132_));
  gate1 g110(new_n132_, new_n129_, 1'b0, 1'b0, 1'b0, new_n95_, new_n133_);
  gate1 g111(n, l, 1'b1, 1'b1, 1'b1, 1'b0, new_n134_);
  gate1 g112(new_n134_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n135_);
  gate1 g113(new_n25_, j, 1'b0, 1'b0, 1'b0, new_n35_, new_n136_);
  gate1 g114(new_n136_, new_n135_, 1'b0, 1'b1, 1'b1, 1'b1, new_n137_);
  gate1 g115(new_n137_, new_n90_, 1'b0, 1'b0, 1'b0, new_n130_, new_n138_);
  gate1 g116(new_n68_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n139_);
  gate1 g117(new_n94_, new_n90_, 1'b0, 1'b0, 1'b0, new_n139_, new_n140_);
  gate1 g118(new_n137_, new_n91_, 1'b0, 1'b0, 1'b0, new_n96_, new_n141_);
  gate1 g119(new_n141_, new_n140_, 1'b0, 1'b0, 1'b0, new_n138_, new_n142_);
  gate1 g120(n, m, 1'b1, 1'b1, 1'b1, 1'b0, new_n143_);
  oai21  g121(.a(new_n142_), .b(new_n133_), .c(new_n143_), .O(new_n144_));
  gate1 g122(m, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n145_);
  gate1 g123(new_n142_, new_n133_, 1'b0, 1'b1, 1'b1, 1'b1, new_n146_);
  gate1 g124(new_n146_, n, 1'b0, 1'b0, 1'b0, new_n145_, new_n147_);
  gate1 g125(new_n67_, ew_n47_), .c(new_n31_, 1'b0, 1'b1, new_n47_, 1'b1, new_n148_);
  gate1 g126(n, new_n23_, 1'b0, 1'b1, 1'b1, 1'b1, new_n149_);
  gate1 g127(new_n149_, new_n53_, 1'b1, 1'b1, 1'b1, 1'b0, new_n150_);
  gate1 g128(new_n52_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n151_);
  gate1 g129(k, i, 1'b0, 1'b1, 1'b1, 1'b1, new_n152_);
  gate1 g130(l, ), .c(new_n152_, 1'b0, 1'b1, k, 1'b1, new_n153_);
  gate1 g131(new_n153_, new_n151_, 1'b0, 1'b1, 1'b1, 1'b1, new_n154_);
  gate1 g132(new_n52_, new_n44_, 1'b0, 1'b0, 1'b0, l, new_n155_);
  gate1 g133(new_n27_, new_n23_, 1'b0, 1'b0, 1'b0, new_n32_, new_n156_);
  oai21  g134(.a(new_n156_), .b(new_n73_), .c(new_n155_), .O(new_n157_));
  gate1 g135(l, new_n35_, 1'b0, 1'b0, 1'b0, 1'b1, new_n158_);
  gate1 g136(new_n149_, new_n32_, 1'b0, 1'b0, 1'b0, new_n31_, new_n159_);
  gate1 g137(new_n27_, j, 1'b0, 1'b0, 1'b0, e, new_n160_);
  oai22  g138(.a(new_n160_), .b(new_n158_), .c(new_n159_), .d(new_n59_), .O(new_n161_));
  gate1 g139(new_n161_, new_n157_, 1'b0, 1'b1, 1'b1, 1'b1, new_n162_);
  gate1 g140(l, new_n25_, 1'b0, 1'b0, 1'b0, i, new_n163_);
  gate1 g141(new_n163_, new_n151_, 1'b0, 1'b1, 1'b1, 1'b1, new_n164_);
  gate1 g142(new_n25_, i, 1'b0, 1'b1, 1'b1, 1'b1, new_n165_);
  oai21  g143(.a(new_n165_), .b(l), .c(new_n149_), .O(new_n166_));
  gate1 g144(new_n166_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n167_);
  aoi22  g145(.a(new_n167_), .b(new_n49_), .c(new_n164_), .d(new_n106_), .O(new_n168_));
  gate1 g146(new_n63_, ew_n25_), .c(n, 1'b0, 1'b1, new_n25_, 1'b1, new_n169_);
  gate1 g147(l, k, 1'b0, 1'b1, 1'b1, 1'b1, new_n170_);
  gate1 g148(n, j, 1'b0, 1'b0, 1'b0, i, new_n171_);
  gate1 g149(new_n171_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n172_);
  gate1 g150(k, new_n23_, 1'b0, 1'b0, 1'b0, 1'b1, new_n173_);
  gate1 g151(new_n173_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n174_);
  gate1 g152(new_n27_, l, 1'b0, 1'b0, 1'b0, new_n35_, new_n175_);
  gate1 g153(new_n175_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n176_);
  aoi22  g154(.a(new_n176_), .b(new_n174_), .c(new_n172_), .d(new_n170_), .O(new_n177_));
  gate1 g155(new_n177_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n178_);
  gate1 g156(new_n169_, ew_n100_), .c(new_n178_, 1'b0, 1'b1, new_n100_, 1'b1, new_n179_);
  gate1 g157(new_n179_, new_n168_, 1'b0, 1'b0, 1'b0, new_n162_, new_n180_);
  gate1 g158(new_n154_, ew_n68_), .c(new_n180_, 1'b0, 1'b1, new_n68_, 1'b1, new_n181_);
  gate1 g159(new_n170_, ), .c(new_n165_, 1'b0, 1'b1, i, 1'b1, new_n182_);
  gate1 g160(new_n182_, new_n151_, 1'b0, 1'b1, 1'b1, 1'b1, new_n183_);
  gate1 g161(new_n183_, new_n67_, 1'b0, 1'b0, 1'b0, new_n47_, new_n184_);
  gate1 g162(new_n36_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n185_);
  gate1 g163(new_n68_, new_n185_, 1'b0, 1'b0, 1'b0, e, new_n186_);
  gate1 g164(new_n186_, new_n184_, 1'b0, 1'b0, 1'b0, new_n181_, new_n187_);
  gate1 g165(new_n150_, ew_n148_), .c(new_n187_, 1'b0, 1'b1, new_n148_, 1'b1, new_n188_);
  gate1 g166(new_n188_, new_n147_, 1'b0, 1'b0, 1'b0, new_n144_, o);
  gate1 g167(f, b, 1'b0, 1'b0, 1'b0, 1'b1, new_n190_);
  gate1 g168(new_n190_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n191_);
  gate1 g169(new_n26_, k, 1'b0, 1'b0, 1'b0, new_n23_, new_n192_);
  gate1 g170(new_n192_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n193_);
  gate1 g171(new_n193_, n, 1'b0, 1'b0, 1'b0, 1'b1, new_n194_);
  gate1 g172(new_n194_, new_n65_, 1'b0, 1'b0, 1'b0, new_n61_, new_n195_);
  gate1 g173(new_n195_, new_n191_, 1'b0, 1'b0, 1'b0, 1'b1, new_n196_);
  gate1 g174(f, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n197_);
  gate1 g175(new_n58_, new_n197_, 1'b1, 1'b1, 1'b1, 1'b0, new_n198_);
  gate1 g176(new_n198_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n199_);
  gate1 g177(e, ew_n31_), .c(new_n23_, 1'b0, 1'b1, new_n31_, 1'b1, new_n200_);
  gate1 g178(n, new_n35_, 1'b0, 1'b0, 1'b0, 1'b1, new_n201_);
  gate1 g179(b, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n202_);
  gate1 g180(f, new_n202_, 1'b0, 1'b0, 1'b0, 1'b1, new_n203_);
  gate1 g181(new_n203_, new_n201_, new_n41_, 1'b1, 1'b1, 1'b1, new_n204_);
  gate1 g182(new_n204_, new_n200_, 1'b0, 1'b0, 1'b0, 1'b1, new_n205_);
  gate1 g183(new_n197_, b, 1'b0, 1'b0, 1'b0, 1'b1, new_n206_);
  gate1 g184(new_n206_, new_n201_, 1'b0, 1'b1, 1'b1, 1'b1, new_n207_);
  gate1 g185(new_n197_, new_n202_, 1'b0, 1'b0, 1'b0, 1'b1, new_n208_);
  gate1 g186(new_n208_, new_n42_, 1'b0, 1'b1, 1'b1, 1'b1, new_n209_);
  aoi22  g187(.a(new_n209_), .b(new_n40_), .c(new_n207_), .d(new_n200_), .O(new_n210_));
  gate1 g188(new_n201_, new_n42_, 1'b0, 1'b1, 1'b1, 1'b1, new_n211_);
  gate1 g189(new_n190_, new_n41_, 1'b0, 1'b1, 1'b1, 1'b1, new_n212_);
  gate1 g190(new_n201_, new_n173_, 1'b0, 1'b1, 1'b1, 1'b1, new_n213_);
  aoi22  g191(.a(new_n213_), .b(new_n100_), .c(new_n212_), .d(new_n211_), .O(new_n214_));
  gate1 g192(new_n214_, new_n210_, 1'b0, 1'b0, 1'b0, new_n205_, new_n215_);
  gate1 g193(new_n37_, new_n202_, 1'b0, 1'b0, 1'b0, 1'b1, new_n216_);
  gate1 g194(new_n208_, new_n30_, 1'b0, 1'b0, 1'b0, 1'b1, new_n217_);
  gate1 g195(new_n217_, new_n216_, 1'b0, 1'b0, 1'b0, 1'b1, new_n218_);
  gate1 g196(new_n218_, new_n215_, 1'b0, 1'b1, 1'b1, 1'b1, new_n219_);
  gate1 g197(new_n219_, new_n199_, 1'b0, 1'b0, 1'b0, new_n196_, new_n220_);
  gate1 g198(j, i, 1'b0, 1'b0, 1'b0, b, new_n221_);
  gate1 g199(new_n221_, new_n75_, 1'b0, 1'b1, 1'b1, 1'b1, new_n222_);
  gate1 g200(new_n191_, new_n23_, 1'b0, 1'b0, 1'b0, i, new_n223_);
  oai22  g201(.a(new_n223_), .b(new_n75_), .c(new_n70_), .d(new_n202_), .O(new_n224_));
  gate1 g202(new_n222_, ew_n220_), .c(new_n224_, 1'b0, 1'b1, new_n220_, 1'b1, new_n225_);
  gate1 g203(new_n218_, new_n215_, new_n198_, 1'b1, 1'b1, 1'b1, new_n226_);
  gate1 g204(new_n226_, new_n196_, 1'b0, 1'b0, 1'b0, new_n82_, new_n227_);
  gate1 g205(new_n220_, new_n71_, 1'b0, 1'b0, 1'b0, 1'b1, new_n228_);
  gate1 g206(new_n228_, new_n227_, 1'b0, 1'b0, 1'b0, new_n225_, new_n229_);
  gate1 g207(new_n96_, a, 1'b0, 1'b0, 1'b0, 1'b1, new_n230_);
  gate1 g208(new_n230_, new_n229_, 1'b1, 1'b0, 1'b0, 1'b0, new_n231_);
  gate1 g209(new_n231_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n232_);
  gate1 g210(k, new_n35_, 1'b0, 1'b0, 1'b0, new_n202_, new_n233_);
  gate1 g211(new_n233_, new_n93_, 1'b0, 1'b1, 1'b1, 1'b1, new_n234_);
  gate1 g212(new_n234_, new_n232_, 1'b0, 1'b0, 1'b0, 1'b1, new_n235_);
  aoi22  g213(.a(new_n89_), .b(new_n72_), .c(new_n88_), .d(new_n77_), .O(new_n236_));
  gate1 g214(new_n74_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n237_);
  gate1 g215(new_n191_, new_n71_, 1'b0, 1'b0, 1'b0, new_n25_, new_n238_);
  oai21  g216(.a(new_n229_), .b(new_n237_), .c(new_n238_), .O(new_n239_));
  gate1 g217(n, new_n25_, 1'b0, 1'b0, 1'b0, j, new_n240_);
  gate1 g218(new_n240_, new_n158_, 1'b0, 1'b1, 1'b1, 1'b1, new_n241_);
  gate1 g219(new_n241_, new_n229_, 1'b1, 1'b1, 1'b1, 1'b0, new_n242_);
  gate1 g220(new_n242_, new_n239_, 1'b0, 1'b0, 1'b0, new_n236_, new_n243_);
  gate1 g221(new_n93_, i, new_n202_, 1'b1, 1'b1, 1'b1, new_n244_);
  gate1 g222(new_n244_, new_n231_, 1'b0, 1'b0, 1'b0, 1'b1, new_n245_);
  gate1 g223(new_n245_, new_n243_, 1'b0, 1'b0, 1'b0, new_n235_, new_n246_);
  gate1 g224(new_n246_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n247_);
  gate1 g225(new_n89_, ew_n72_), .c(new_n139_, 1'b0, 1'b1, new_n72_, 1'b1, new_n248_);
  gate1 g226(new_n220_, new_n94_, 1'b1, 1'b1, 1'b1, 1'b0, new_n249_);
  gate1 g227(new_n249_, new_n248_, 1'b0, 1'b0, 1'b0, new_n239_, new_n250_);
  gate1 g228(new_n239_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n251_);
  gate1 g229(new_n242_, new_n251_, 1'b0, 1'b0, 1'b0, 1'b1, new_n252_);
  oai21  g230(.a(new_n252_), .b(new_n236_), .c(new_n250_), .O(new_n253_));
  gate1 g231(new_n241_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n254_);
  gate1 g232(new_n254_, new_n229_, 1'b0, 1'b1, 1'b1, 1'b1, new_n255_);
  gate1 g233(new_n255_, new_n239_, 1'b0, 1'b0, 1'b0, 1'b1, new_n256_);
  gate1 g234(new_n255_, new_n251_, 1'b0, 1'b0, 1'b0, new_n236_, new_n257_);
  oai21  g235(.a(new_n256_), .b(new_n236_), .c(new_n257_), .O(new_n258_));
  gate1 g236(new_n258_, new_n253_, 1'b0, 1'b1, 1'b1, 1'b1, new_n259_);
  gate1 g237(new_n248_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n260_);
  gate1 g238(new_n249_, new_n260_, 1'b0, 1'b0, 1'b0, new_n251_, new_n261_);
  gate1 g239(new_n109_, new_n27_, l, 1'b1, 1'b1, 1'b1, new_n262_);
  gate1 g240(new_n229_, new_n96_, 1'b0, 1'b1, 1'b1, 1'b1, new_n263_);
  gate1 g241(new_n262_, new_n229_, 1'b0, 1'b0, 1'b0, new_n96_, new_n264_);
  gate1 g242(l, k, 1'b1, 1'b1, 1'b1, 1'b0, new_n265_);
  gate1 g243(new_n265_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n266_);
  oai22  g244(.a(new_n266_), .b(new_n56_), .c(new_n63_), .d(new_n26_), .O(new_n267_));
  gate1 g245(new_n267_, n, 1'b0, 1'b0, 1'b0, new_n202_, new_n268_);
  gate1 g246(new_n268_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n269_);
  gate1 g247(new_n269_, new_n68_, 1'b0, 1'b0, 1'b0, a, new_n270_);
  gate1 g248(new_n220_, n, 1'b0, 1'b0, 1'b0, 1'b1, new_n271_);
  gate1 g249(new_n123_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n272_);
  gate1 g250(new_n26_, j, 1'b0, 1'b0, 1'b0, new_n35_, new_n273_);
  gate1 g251(new_n273_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n274_);
  gate1 g252(new_n272_, ), .c(new_n274_, 1'b0, 1'b1, l, 1'b1, new_n275_);
  gate1 g253(new_n275_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n276_);
  oai21  g254(.a(new_n80_), .b(new_n46_), .c(new_n276_), .O(new_n277_));
  oai22  g255(.a(new_n277_), .b(new_n271_), .c(new_n270_), .d(new_n220_), .O(new_n278_));
  gate1 g256(new_n136_, l, 1'b0, 1'b1, 1'b1, 1'b1, new_n279_);
  gate1 g257(new_n279_, new_n220_, 1'b0, 1'b0, 1'b0, n, new_n280_);
  gate1 g258(new_n226_, new_n196_, 1'b0, 1'b0, 1'b0, new_n139_, new_n281_);
  oai21  g259(.a(new_n281_), .b(new_n125_), .c(new_n280_), .O(new_n282_));
  gate1 g260(new_n282_, new_n278_, 1'b0, 1'b1, 1'b1, 1'b1, new_n283_);
  oai21  g261(.a(new_n80_), .b(new_n46_), .c(a), .O(new_n284_));
  gate1 g262(new_n267_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n285_);
  oai21  g263(.a(new_n63_), .b(k), .c(new_n285_), .O(new_n286_));
  gate1 g264(n, b, 1'b1, 1'b1, 1'b1, 1'b0, new_n287_);
  gate1 g265(new_n287_, new_n286_, 1'b0, 1'b0, 1'b0, new_n284_, new_n288_);
  gate1 g266(new_n104_, new_n103_, 1'b0, 1'b0, 1'b0, f, new_n289_);
  gate1 g267(new_n109_, new_n27_, 1'b0, 1'b1, 1'b1, 1'b1, new_n290_);
  gate1 g268(new_n290_, new_n100_, 1'b0, 1'b0, 1'b0, b, new_n291_);
  gate1 g269(b, a, 1'b0, 1'b1, 1'b1, 1'b1, new_n292_);
  gate1 g270(new_n292_, new_n290_, 1'b0, 1'b0, 1'b0, l, new_n293_);
  gate1 g271(new_n293_, new_n291_, 1'b0, 1'b0, 1'b0, new_n289_, new_n294_);
  gate1 g272(new_n25_, new_n23_, 1'b0, 1'b0, 1'b0, i, new_n295_);
  gate1 g273(new_n295_, new_n27_, 1'b0, 1'b1, 1'b1, 1'b1, new_n296_);
  gate1 g274(new_n208_, new_n48_, 1'b0, 1'b1, 1'b1, 1'b1, new_n297_);
  gate1 g275(new_n297_, new_n296_, 1'b0, 1'b0, 1'b0, l, new_n298_);
  gate1 g276(new_n48_, new_n197_, 1'b0, 1'b0, 1'b0, b, new_n299_);
  gate1 g277(new_n299_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n300_);
  gate1 g278(new_n55_, new_n26_, 1'b0, 1'b0, 1'b0, new_n25_, new_n301_);
  gate1 g279(new_n301_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n302_);
  aoi22  g280(.a(new_n302_), .b(new_n287_), .c(new_n300_), .d(new_n296_), .O(new_n303_));
  gate1 g281(new_n190_, new_n48_, 1'b0, 1'b1, 1'b1, 1'b1, new_n304_);
  gate1 g282(new_n48_, f, 1'b0, 1'b0, 1'b0, new_n202_, new_n305_);
  gate1 g283(new_n305_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n306_);
  oai21  g284(.a(new_n306_), .b(new_n304_), .c(new_n296_), .O(new_n307_));
  gate1 g285(new_n307_, new_n303_, 1'b0, 1'b0, 1'b0, new_n298_, new_n308_);
  gate1 g286(new_n308_, new_n294_, 1'b0, 1'b1, 1'b1, 1'b1, new_n309_);
  oai21  g287(.a(new_n288_), .b(new_n220_), .c(new_n309_), .O(new_n310_));
  gate1 g288(new_n286_, new_n148_, 1'b0, 1'b0, 1'b0, b, new_n311_);
  gate1 g289(new_n269_, new_n220_, 1'b0, 1'b0, 1'b0, new_n284_, new_n312_);
  oai21  g290(.a(new_n311_), .b(new_n271_), .c(new_n312_), .O(new_n313_));
  gate1 g291(new_n313_, new_n310_, 1'b0, 1'b1, 1'b1, 1'b1, new_n314_);
  gate1 g292(new_n314_, new_n283_, 1'b0, 1'b0, 1'b0, new_n264_, new_n315_);
  gate1 g293(new_n263_, ew_n262_), .c(new_n315_, 1'b0, 1'b1, new_n262_, 1'b1, new_n316_);
  gate1 g294(new_n316_, new_n261_, 1'b0, 1'b0, 1'b0, 1'b1, new_n317_);
  gate1 g295(new_n220_, new_n93_, new_n92_, 1'b1, 1'b1, 1'b1, new_n318_);
  gate1 g296(new_n318_, new_n248_, 1'b0, 1'b0, 1'b0, new_n251_, new_n319_);
  gate1 g297(new_n318_, new_n260_, 1'b0, 1'b0, 1'b0, new_n239_, new_n320_);
  gate1 g298(new_n320_, new_n319_, 1'b0, 1'b0, 1'b0, 1'b1, new_n321_);
  gate1 g299(new_n321_, new_n317_, 1'b0, 1'b1, 1'b1, 1'b1, new_n322_);
  gate1 g300(new_n322_, new_n259_, 1'b0, 1'b0, 1'b0, new_n247_, new_n323_);
  gate1 g301(new_n146_, m, 1'b0, 1'b1, 1'b1, 1'b1, new_n324_);
  gate1 g302(new_n324_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n325_);
  gate1 g303(new_n325_, new_n323_, 1'b0, 1'b0, 1'b0, n, new_n326_);
  gate1 g304(new_n323_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n327_);
  gate1 g305(new_n324_, new_n327_, 1'b0, 1'b0, 1'b0, n, new_n328_);
  gate1 g306(new_n220_, new_n185_, 1'b0, 1'b0, 1'b0, f, new_n329_);
  gate1 g307(new_n226_, new_n196_, 1'b0, 1'b0, 1'b0, new_n183_, new_n330_);
  gate1 g308(l, b, 1'b1, 1'b1, 1'b1, 1'b0, new_n331_);
  gate1 g309(new_n331_, new_n169_, 1'b0, 1'b0, 1'b0, 1'b1, new_n332_);
  gate1 g310(new_n197_, b, 1'b0, 1'b1, 1'b1, 1'b1, new_n333_);
  gate1 g311(f, b, 1'b0, 1'b1, 1'b1, 1'b1, new_n334_);
  gate1 g312(new_n59_, n, new_n23_, 1'b1, 1'b1, 1'b1, new_n335_);
  aoi22  g313(.a(new_n335_), .b(new_n334_), .c(new_n333_), .d(new_n164_), .O(new_n336_));
  gate1 g314(new_n336_, new_n332_, 1'b0, 1'b0, 1'b0, 1'b1, new_n337_);
  gate1 g315(new_n41_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n338_);
  gate1 g316(n, j, f, 1'b1, 1'b1, 1'b1, new_n339_);
  gate1 g317(new_n339_, new_n338_, 1'b0, 1'b0, 1'b0, i, new_n340_);
  gate1 g318(new_n176_, j, 1'b0, 1'b0, 1'b0, f, new_n341_);
  gate1 g319(f, new_n202_, 1'b0, 1'b1, 1'b1, 1'b1, new_n342_);
  gate1 g320(new_n342_, new_n52_, 1'b0, 1'b0, 1'b0, l, new_n343_);
  gate1 g321(new_n343_, new_n341_, 1'b0, 1'b0, 1'b0, new_n340_, new_n344_);
  oai21  g322(.a(new_n190_), .b(new_n166_), .c(new_n177_), .O(new_n345_));
  gate1 g323(new_n345_, new_n344_, new_n337_, 1'b1, 1'b1, 1'b1, new_n346_);
  gate1 g324(new_n346_, new_n330_, 1'b0, 1'b0, 1'b0, new_n329_, new_n347_);
  gate1 g325(new_n220_, new_n27_, 1'b0, 1'b0, 1'b0, 1'b1, new_n348_);
  gate1 g326(new_n53_, j, 1'b0, 1'b0, 1'b0, b, new_n349_);
  oai21  g327(.a(new_n265_), .b(new_n152_), .c(new_n23_), .O(new_n350_));
  gate1 g328(new_n350_, ew_n349_), .c(new_n348_, 1'b0, 1'b1, new_n349_, 1'b1, new_n351_);
  gate1 g329(new_n351_, new_n347_, 1'b0, 1'b1, 1'b1, 1'b1, new_n352_);
  gate1 g330(new_n352_, new_n328_, 1'b0, 1'b0, 1'b0, new_n326_, p);
  gate1 g331(new_n229_, new_n90_, 1'b0, 1'b0, 1'b0, new_n96_, new_n354_);
  gate1 g332(new_n239_, new_n90_, 1'b0, 1'b0, 1'b0, new_n96_, new_n355_);
  gate1 g333(new_n239_, new_n229_, 1'b0, 1'b0, 1'b0, 1'b1, new_n356_);
  gate1 g334(new_n356_, new_n355_, 1'b0, 1'b0, 1'b0, new_n354_, new_n357_);
  gate1 g335(g, c, 1'b1, 1'b1, 1'b1, 1'b0, new_n358_);
  gate1 g336(new_n358_, new_n195_, 1'b0, 1'b0, 1'b0, 1'b1, new_n359_);
  gate1 g337(g, c, 1'b0, 1'b1, 1'b1, 1'b1, new_n360_);
  gate1 g338(new_n360_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n361_);
  gate1 g339(c, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n362_);
  gate1 g340(new_n37_, new_n362_, 1'b0, 1'b0, 1'b0, 1'b1, new_n363_);
  gate1 g341(new_n206_, ew_n106_), .c(new_n333_, 1'b0, 1'b1, new_n106_, 1'b1, new_n364_);
  gate1 g342(g, new_n362_, 1'b0, 1'b0, 1'b0, 1'b1, new_n365_);
  gate1 g343(new_n365_, new_n39_, new_n41_, 1'b1, 1'b1, 1'b1, new_n366_);
  gate1 g344(new_n366_, new_n364_, 1'b0, 1'b0, 1'b0, 1'b1, new_n367_);
  gate1 g345(new_n331_, new_n213_, 1'b0, 1'b0, 1'b0, 1'b1, new_n368_);
  gate1 g346(new_n368_, new_n367_, 1'b0, 1'b0, 1'b0, new_n363_, new_n369_);
  gate1 g347(new_n361_, ew_n30_), .c(new_n369_, 1'b0, 1'b1, new_n30_, 1'b1, new_n370_);
  gate1 g348(g, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n371_);
  oai21  g349(.a(new_n342_), .b(new_n42_), .c(new_n203_), .O(new_n372_));
  gate1 g350(new_n201_, new_n41_, 1'b0, 1'b1, 1'b1, 1'b1, new_n373_);
  gate1 g351(new_n373_, new_n372_, 1'b0, 1'b0, 1'b0, new_n358_, new_n374_);
  gate1 g352(new_n371_, c, 1'b0, 1'b0, 1'b0, 1'b1, new_n375_);
  gate1 g353(new_n375_, new_n39_, 1'b0, 1'b1, 1'b1, 1'b1, new_n376_);
  gate1 g354(new_n376_, new_n364_, 1'b0, 1'b0, 1'b0, 1'b1, new_n377_);
  gate1 g355(new_n372_, new_n360_, 1'b0, 1'b0, 1'b0, new_n40_, new_n378_);
  gate1 g356(new_n378_, new_n377_, 1'b0, 1'b0, 1'b0, new_n374_, new_n379_);
  gate1 g357(new_n58_, ew_n371_), .c(new_n379_, 1'b0, 1'b1, new_n371_, 1'b1, new_n380_);
  gate1 g358(new_n380_, new_n370_, 1'b0, 1'b0, 1'b0, new_n359_, new_n381_);
  gate1 g359(j, i, 1'b0, 1'b0, 1'b0, c, new_n382_);
  gate1 g360(new_n382_, new_n75_, 1'b0, 1'b1, 1'b1, 1'b1, new_n383_);
  gate1 g361(new_n358_, new_n23_, 1'b0, 1'b0, 1'b0, i, new_n384_);
  oai22  g362(.a(new_n384_), .b(new_n75_), .c(new_n70_), .d(new_n362_), .O(new_n385_));
  gate1 g363(new_n383_, ew_n381_), .c(new_n385_, 1'b0, 1'b1, new_n381_, 1'b1, new_n386_);
  gate1 g364(new_n361_, new_n30_, 1'b0, 1'b0, 1'b0, 1'b1, new_n387_);
  aoi22  g365(.a(new_n366_), .b(new_n364_), .c(new_n331_), .d(new_n213_), .O(new_n388_));
  gate1 g366(new_n388_, new_n363_, 1'b0, 1'b0, 1'b0, new_n387_, new_n389_);
  gate1 g367(new_n58_, new_n371_, 1'b0, 1'b0, 1'b0, 1'b1, new_n390_);
  gate1 g368(new_n379_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n391_);
  gate1 g369(new_n391_, new_n390_, 1'b0, 1'b0, 1'b0, 1'b1, new_n392_);
  gate1 g370(new_n392_, new_n389_, 1'b0, 1'b1, 1'b1, 1'b1, new_n393_);
  gate1 g371(new_n393_, new_n359_, 1'b0, 1'b0, 1'b0, new_n82_, new_n394_);
  gate1 g372(new_n381_, new_n71_, 1'b0, 1'b0, 1'b0, 1'b1, new_n395_);
  gate1 g373(new_n395_, new_n394_, 1'b0, 1'b0, 1'b0, new_n386_, new_n396_);
  gate1 g374(new_n358_, new_n71_, 1'b0, 1'b0, 1'b0, new_n25_, new_n397_);
  oai21  g375(.a(new_n396_), .b(new_n237_), .c(new_n397_), .O(new_n398_));
  gate1 g376(new_n398_, new_n241_, 1'b1, 1'b1, 1'b1, 1'b0, new_n399_);
  gate1 g377(new_n399_, new_n396_, 1'b0, 1'b0, 1'b0, new_n357_, new_n400_);
  gate1 g378(new_n357_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n401_);
  gate1 g379(new_n398_, new_n254_, 1'b0, 1'b1, 1'b1, 1'b1, new_n402_);
  gate1 g380(new_n402_, new_n396_, 1'b0, 1'b0, 1'b0, new_n401_, new_n403_);
  gate1 g381(new_n396_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n404_);
  gate1 g382(new_n402_, new_n404_, 1'b0, 1'b0, 1'b0, new_n357_, new_n405_);
  gate1 g383(new_n405_, new_n403_, 1'b0, 1'b0, 1'b0, new_n400_, new_n406_);
  gate1 g384(new_n406_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n407_);
  gate1 g385(new_n229_, new_n96_, 1'b0, 1'b0, 1'b0, a, new_n408_);
  gate1 g386(new_n96_, b, 1'b0, 1'b0, 1'b0, a, new_n409_);
  gate1 g387(new_n229_, b, 1'b0, 1'b0, 1'b0, 1'b1, new_n410_);
  gate1 g388(new_n410_, new_n409_, 1'b0, 1'b0, 1'b0, new_n408_, new_n411_);
  gate1 g389(new_n411_, new_n396_, 1'b1, 1'b0, 1'b0, 1'b0, new_n412_);
  gate1 g390(k, new_n35_, 1'b0, 1'b0, 1'b0, new_n362_, new_n413_);
  gate1 g391(new_n413_, new_n93_, 1'b0, 1'b1, 1'b1, 1'b1, new_n414_);
  gate1 g392(new_n414_, new_n412_, 1'b0, 1'b0, 1'b0, 1'b1, new_n415_);
  gate1 g393(new_n404_, new_n263_, 1'b0, 1'b0, 1'b0, new_n262_, new_n416_);
  gate1 g394(new_n220_, new_n68_, 1'b0, 1'b0, 1'b0, a, new_n417_);
  oai21  g395(.a(new_n220_), .b(new_n148_), .c(b), .O(new_n418_));
  gate1 g396(new_n418_, new_n417_, 1'b0, 1'b0, 1'b0, 1'b1, new_n419_);
  gate1 g397(new_n267_, new_n362_, 1'b1, 1'b1, 1'b1, 1'b0, new_n420_);
  gate1 g398(new_n420_, new_n381_, 1'b0, 1'b0, 1'b0, n, new_n421_);
  gate1 g399(new_n421_, new_n419_, 1'b0, 1'b1, 1'b1, 1'b1, new_n422_);
  gate1 g400(new_n267_, new_n362_, 1'b0, 1'b0, 1'b0, 1'b1, new_n423_);
  gate1 g401(new_n423_, new_n381_, new_n27_, 1'b1, 1'b1, 1'b1, new_n424_);
  gate1 g402(new_n424_, ew_n419_), .c(new_n422_, 1'b0, 1'b1, new_n419_, 1'b1, new_n425_);
  gate1 g403(new_n381_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n426_);
  gate1 g404(new_n286_, c, 1'b1, 1'b1, 1'b1, 1'b0, new_n427_);
  gate1 g405(new_n427_, new_n426_, 1'b0, 1'b0, 1'b0, n, new_n428_);
  gate1 g406(new_n428_, new_n419_, 1'b1, 1'b0, 1'b0, 1'b0, new_n429_);
  gate1 g407(new_n393_, ew_n359_), .c(new_n27_, 1'b0, 1'b1, new_n359_, 1'b1, new_n430_);
  gate1 g408(new_n427_, new_n430_, 1'b0, 1'b0, 1'b0, new_n419_, new_n431_);
  gate1 g409(new_n431_, new_n429_, 1'b0, 1'b0, 1'b0, new_n425_, new_n432_);
  gate1 g410(new_n229_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n433_);
  gate1 g411(new_n433_, new_n130_, 1'b0, 1'b0, 1'b0, 1'b1, new_n434_);
  gate1 g412(new_n396_, new_n434_, 1'b0, 1'b0, 1'b0, new_n262_, new_n435_);
  gate1 g413(new_n125_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n436_);
  gate1 g414(new_n220_, new_n68_, 1'b0, 1'b1, 1'b1, 1'b1, new_n437_);
  gate1 g415(new_n426_, new_n437_, 1'b0, 1'b0, 1'b0, new_n436_, new_n438_);
  gate1 g416(new_n430_, new_n281_, 1'b0, 1'b0, 1'b0, new_n276_, new_n439_);
  gate1 g417(new_n381_, new_n279_, 1'b0, 1'b0, 1'b0, n, new_n440_);
  gate1 g418(new_n362_, new_n202_, 1'b0, 1'b0, 1'b0, new_n31_, new_n441_);
  gate1 g419(new_n441_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n442_);
  gate1 g420(new_n442_, new_n290_, 1'b0, 1'b0, 1'b0, l, new_n443_);
  gate1 g421(new_n208_, new_n49_, 1'b0, 1'b0, 1'b0, 1'b1, new_n444_);
  gate1 g422(new_n444_, new_n296_, 1'b0, 1'b0, 1'b0, new_n190_, new_n445_);
  gate1 g423(new_n445_, new_n365_, 1'b1, 1'b0, 1'b0, 1'b0, new_n446_);
  oai21  g424(.a(new_n334_), .b(new_n48_), .c(new_n190_), .O(new_n447_));
  gate1 g425(new_n447_, new_n358_, 1'b0, 1'b0, 1'b0, new_n296_, new_n448_);
  gate1 g426(new_n448_, new_n446_, 1'b0, 1'b0, 1'b0, new_n443_, new_n449_);
  gate1 g427(new_n104_, new_n103_, 1'b0, 1'b0, 1'b0, g, new_n450_);
  gate1 g428(new_n292_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n451_);
  gate1 g429(l, c, 1'b1, 1'b1, 1'b1, 1'b0, new_n452_);
  gate1 g430(new_n452_, new_n451_, 1'b0, 1'b0, 1'b0, new_n290_, new_n453_);
  gate1 g431(new_n302_, n, 1'b0, 1'b0, 1'b0, c, new_n454_);
  gate1 g432(new_n454_, new_n453_, 1'b0, 1'b0, 1'b0, new_n450_, new_n455_);
  gate1 g433(new_n295_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n456_);
  gate1 g434(new_n447_, new_n456_, 1'b0, 1'b0, 1'b0, n, new_n457_);
  gate1 g435(l, new_n371_, 1'b0, 1'b0, 1'b0, new_n362_, new_n458_);
  oai22  g436(.a(new_n458_), .b(new_n457_), .c(new_n445_), .d(new_n375_), .O(new_n459_));
  gate1 g437(new_n459_, new_n455_, new_n449_, 1'b1, 1'b1, 1'b1, new_n460_);
  gate1 g438(new_n460_, new_n440_, 1'b1, 1'b1, 1'b1, 1'b0, new_n461_);
  gate1 g439(new_n461_, new_n439_, 1'b1, 1'b1, 1'b1, 1'b0, new_n462_);
  gate1 g440(new_n462_, new_n438_, 1'b0, 1'b0, 1'b0, new_n435_, new_n463_);
  gate1 g441(new_n463_, new_n432_, 1'b0, 1'b1, 1'b1, 1'b1, new_n464_);
  gate1 g442(new_n464_, new_n416_, 1'b0, 1'b0, 1'b0, new_n415_, new_n465_);
  gate1 g443(new_n465_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n466_);
  gate1 g444(new_n103_, new_n35_, 1'b0, 1'b0, 1'b0, c, new_n467_);
  gate1 g445(new_n220_, new_n90_, 1'b0, 1'b0, 1'b0, new_n68_, new_n468_);
  gate1 g446(new_n239_, new_n90_, 1'b0, 1'b0, 1'b0, new_n68_, new_n469_);
  gate1 g447(new_n239_, new_n220_, 1'b0, 1'b0, 1'b0, 1'b1, new_n470_);
  gate1 g448(new_n470_, new_n469_, 1'b0, 1'b0, 1'b0, new_n468_, new_n471_);
  gate1 g449(new_n398_, new_n381_, 1'b1, 1'b0, 1'b0, 1'b0, new_n472_);
  gate1 g450(new_n472_, new_n94_, 1'b0, 1'b0, 1'b0, 1'b1, new_n473_);
  oai22  g451(.a(new_n473_), .b(new_n471_), .c(new_n467_), .d(new_n412_), .O(new_n474_));
  gate1 g452(new_n398_, new_n426_, 1'b1, 1'b0, 1'b0, 1'b0, new_n475_);
  gate1 g453(new_n475_, new_n471_, 1'b0, 1'b0, 1'b0, new_n94_, new_n476_);
  gate1 g454(new_n398_, new_n404_, 1'b0, 1'b0, 1'b0, new_n241_, new_n477_);
  oai21  g455(.a(new_n477_), .b(new_n357_), .c(new_n476_), .O(new_n478_));
  gate1 g456(new_n478_, new_n474_, 1'b0, 1'b1, 1'b1, 1'b1, new_n479_);
  gate1 g457(new_n479_, new_n466_, 1'b0, 1'b0, 1'b0, new_n407_, new_n480_);
  gate1 g458(new_n324_, new_n323_, 1'b0, 1'b0, 1'b0, 1'b1, new_n481_);
  gate1 g459(new_n481_, new_n480_, 1'b0, 1'b0, 1'b0, n, new_n482_);
  gate1 g460(new_n324_, new_n323_, 1'b0, 1'b0, 1'b0, n, new_n483_);
  gate1 g461(new_n483_, new_n480_, 1'b1, 1'b0, 1'b0, 1'b0, new_n484_);
  gate1 g462(new_n381_, new_n185_, 1'b0, 1'b0, 1'b0, g, new_n485_);
  gate1 g463(n, j, g, 1'b1, 1'b1, 1'b1, new_n486_);
  gate1 g464(new_n360_, new_n27_, 1'b0, 1'b0, 1'b0, j, new_n487_);
  gate1 g465(n, new_n371_, 1'b0, 1'b1, 1'b1, 1'b1, new_n488_);
  gate1 g466(new_n488_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n489_);
  gate1 g467(l, j, 1'b0, 1'b0, 1'b0, new_n35_, new_n490_);
  oai22  g468(.a(new_n490_), .b(new_n489_), .c(new_n487_), .d(new_n59_), .O(new_n491_));
  gate1 g469(new_n486_, ew_n452_), .c(new_n491_, 1'b0, 1'b1, new_n452_, 1'b1, new_n492_);
  gate1 g470(new_n486_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n493_);
  gate1 g471(new_n488_, new_n23_, 1'b0, 1'b0, 1'b0, new_n362_, new_n494_);
  oai22  g472(.a(new_n494_), .b(new_n163_), .c(new_n493_), .d(new_n73_), .O(new_n495_));
  gate1 g473(new_n495_, new_n178_, 1'b0, 1'b1, 1'b1, 1'b1, new_n496_);
  aoi22  g474(.a(new_n452_), .b(new_n169_), .c(new_n358_), .d(new_n167_), .O(new_n497_));
  gate1 g475(new_n497_, new_n496_, 1'b0, 1'b0, 1'b0, new_n492_, new_n498_);
  gate1 g476(new_n426_, ew_n183_), .c(new_n498_, 1'b0, 1'b1, new_n183_, 1'b1, new_n499_);
  gate1 g477(new_n499_, new_n485_, 1'b0, 1'b0, 1'b0, 1'b1, new_n500_);
  gate1 g478(new_n381_, new_n27_, 1'b0, 1'b0, 1'b0, 1'b1, new_n501_);
  gate1 g479(new_n53_, j, 1'b0, 1'b0, 1'b0, c, new_n502_);
  gate1 g480(new_n502_, ew_n350_), .c(new_n501_, 1'b0, 1'b1, new_n350_, 1'b1, new_n503_);
  gate1 g481(new_n503_, new_n500_, 1'b0, 1'b1, 1'b1, 1'b1, new_n504_);
  gate1 g482(new_n504_, new_n484_, 1'b0, 1'b0, 1'b0, new_n482_, q);
  gate1 g483(new_n396_, new_n357_, 1'b0, 1'b0, 1'b0, 1'b1, new_n506_);
  gate1 g484(new_n398_, new_n357_, 1'b0, 1'b0, 1'b0, 1'b1, new_n507_);
  gate1 g485(new_n398_, new_n396_, 1'b0, 1'b0, 1'b0, 1'b1, new_n508_);
  gate1 g486(new_n508_, new_n507_, 1'b0, 1'b0, 1'b0, new_n506_, new_n509_);
  gate1 g487(h, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n510_);
  oai21  g488(.a(h), .b(d), .c(new_n30_), .O(new_n511_));
  gate1 g489(n, h, 1'b0, 1'b0, 1'b0, d, new_n512_);
  gate1 g490(new_n512_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n513_);
  gate1 g491(new_n513_, new_n193_, 1'b0, 1'b0, 1'b0, 1'b1, new_n514_);
  gate1 g492(new_n452_, new_n213_, 1'b0, 1'b0, 1'b0, 1'b1, new_n515_);
  gate1 g493(h, d, 1'b1, 1'b1, 1'b1, 1'b0, t);
  gate1 g494(t, new_n193_, 1'b0, 1'b0, 1'b0, new_n35_, new_n517_);
  gate1 g495(new_n517_, new_n515_, 1'b0, 1'b0, 1'b0, new_n514_, new_n518_);
  gate1 g496(new_n518_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n519_);
  gate1 g497(i, d, 1'b0, 1'b1, 1'b1, 1'b1, new_n520_);
  gate1 g498(new_n520_, new_n27_, 1'b0, 1'b0, 1'b0, new_n25_, new_n521_);
  gate1 g499(l, ), .c(new_n521_, 1'b0, 1'b1, j, 1'b1, new_n522_);
  gate1 g500(new_n513_, ew_n64_), .c(new_n522_, 1'b0, 1'b1, new_n64_, 1'b1, new_n523_);
  gate1 g501(new_n523_, new_n519_, 1'b0, 1'b0, 1'b0, new_n511_, new_n524_);
  gate1 g502(new_n58_, ew_n510_), .c(new_n524_, 1'b0, 1'b1, new_n510_, 1'b1, new_n525_);
  gate1 g503(new_n364_, new_n371_, 1'b0, 1'b0, 1'b0, 1'b1, new_n526_);
  gate1 g504(new_n364_, c, 1'b0, 1'b0, 1'b0, 1'b1, new_n527_);
  gate1 g505(new_n527_, new_n526_, 1'b0, 1'b0, 1'b0, new_n375_, new_n528_);
  gate1 g506(d, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n529_);
  gate1 g507(h, new_n529_, 1'b0, 1'b0, 1'b0, 1'b1, new_n530_);
  gate1 g508(new_n530_, new_n39_, new_n41_, 1'b1, 1'b1, 1'b1, new_n531_);
  gate1 g509(new_n531_, new_n528_, 1'b0, 1'b0, 1'b0, 1'b1, new_n532_);
  gate1 g510(new_n39_, h, new_n529_, 1'b1, 1'b1, 1'b1, new_n533_);
  gate1 g511(new_n533_, new_n528_, 1'b0, 1'b0, 1'b0, 1'b1, new_n534_);
  gate1 g512(new_n534_, new_n532_, 1'b0, 1'b0, 1'b0, 1'b1, new_n535_);
  gate1 g513(h, d, 1'b0, 1'b1, 1'b1, 1'b1, new_n536_);
  gate1 g514(new_n536_, new_n50_, 1'b0, 1'b0, 1'b0, n, new_n537_);
  gate1 g515(new_n513_, new_n60_, 1'b0, 1'b0, 1'b0, 1'b1, new_n538_);
  gate1 g516(new_n538_, ew_n537_), .c(new_n528_, 1'b0, 1'b1, new_n537_, 1'b1, new_n539_);
  gate1 g517(new_n539_, new_n535_, 1'b0, 1'b1, 1'b1, 1'b1, new_n540_);
  gate1 g518(new_n540_, new_n525_, 1'b0, 1'b0, 1'b0, 1'b1, new_n541_);
  gate1 g519(new_n541_, new_n76_, 1'b0, 1'b0, 1'b0, d, new_n542_);
  gate1 g520(new_n58_, new_n510_, 1'b0, 1'b0, 1'b0, 1'b1, new_n543_);
  gate1 g521(new_n524_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n544_);
  gate1 g522(new_n544_, new_n543_, 1'b0, 1'b0, 1'b0, 1'b1, new_n545_);
  oai21  g523(.a(new_n533_), .b(new_n531_), .c(new_n528_), .O(new_n546_));
  gate1 g524(new_n528_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n547_);
  gate1 g525(new_n547_, new_n536_, 1'b0, 1'b0, 1'b0, new_n40_, new_n548_);
  gate1 g526(new_n547_, new_n513_, 1'b0, 1'b0, 1'b0, new_n60_, new_n549_);
  gate1 g527(new_n549_, new_n548_, 1'b0, 1'b0, 1'b0, new_n546_, new_n550_);
  oai21  g528(.a(new_n550_), .b(new_n545_), .c(new_n71_), .O(new_n551_));
  gate1 g529(new_n550_, new_n545_, 1'b0, 1'b1, 1'b1, 1'b1, new_n552_);
  gate1 g530(t, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n553_);
  gate1 g531(new_n553_, new_n24_, 1'b0, 1'b1, 1'b1, 1'b1, new_n554_);
  aoi22  g532(.a(new_n554_), .b(new_n84_), .c(new_n71_), .d(d), .O(new_n555_));
  gate1 g533(new_n555_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n556_);
  gate1 g534(new_n552_, ew_n82_), .c(new_n556_, 1'b0, 1'b1, new_n82_, 1'b1, new_n557_);
  gate1 g535(new_n557_, new_n551_, 1'b0, 1'b0, 1'b0, new_n542_, new_n558_);
  gate1 g536(t, new_n71_, 1'b0, 1'b0, 1'b0, new_n25_, new_n559_);
  oai21  g537(.a(new_n558_), .b(new_n237_), .c(new_n559_), .O(new_n560_));
  gate1 g538(new_n136_, new_n27_, new_n26_, 1'b1, 1'b1, 1'b1, new_n561_);
  gate1 g539(new_n561_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n562_);
  gate1 g540(new_n562_, new_n560_, new_n558_, 1'b1, 1'b1, 1'b1, new_n563_);
  gate1 g541(new_n561_, new_n560_, 1'b0, 1'b0, 1'b0, new_n558_, new_n564_);
  gate1 g542(new_n564_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n565_);
  oai21  g543(.a(new_n565_), .b(new_n563_), .c(new_n509_), .O(new_n566_));
  gate1 g544(new_n471_, new_n381_, 1'b0, 1'b0, 1'b0, 1'b1, new_n567_);
  oai21  g545(.a(new_n471_), .b(new_n381_), .c(new_n398_), .O(new_n568_));
  gate1 g546(new_n560_, new_n552_, 1'b0, 1'b0, 1'b0, 1'b1, new_n569_);
  gate1 g547(new_n540_, ew_n525_), .c(new_n529_, 1'b0, 1'b1, new_n525_, 1'b1, new_n570_);
  gate1 g548(new_n540_, new_n525_, 1'b0, 1'b0, 1'b0, new_n82_, new_n571_);
  gate1 g549(new_n555_, new_n571_, 1'b0, 1'b0, 1'b0, new_n551_, new_n572_);
  gate1 g550(new_n570_, ew_n76_), .c(new_n572_, 1'b0, 1'b1, new_n76_, 1'b1, new_n573_);
  gate1 g551(new_n573_, new_n74_, 1'b0, 1'b0, 1'b0, 1'b1, new_n574_);
  gate1 g552(new_n574_, new_n559_, 1'b0, 1'b0, 1'b0, new_n541_, new_n575_);
  gate1 g553(new_n192_, new_n27_, new_n35_, 1'b1, 1'b1, 1'b1, new_n576_);
  gate1 g554(new_n576_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n577_);
  gate1 g555(new_n575_, ew_n569_), .c(new_n577_, 1'b0, 1'b1, new_n569_, 1'b1, new_n578_);
  gate1 g556(new_n578_, new_n568_, 1'b0, 1'b0, 1'b0, new_n567_, new_n579_);
  gate1 g557(new_n568_, new_n567_, 1'b0, 1'b0, 1'b0, 1'b1, new_n580_);
  gate1 g558(new_n576_, new_n575_, 1'b0, 1'b0, 1'b0, new_n569_, new_n581_);
  gate1 g559(new_n581_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n582_);
  gate1 g560(new_n582_, new_n580_, 1'b0, 1'b0, 1'b0, 1'b1, new_n583_);
  gate1 g561(new_n583_, new_n579_, 1'b0, 1'b0, 1'b0, new_n566_, new_n584_);
  gate1 g562(new_n584_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n585_);
  gate1 g563(new_n411_, new_n396_, 1'b0, 1'b0, 1'b0, 1'b1, new_n586_);
  oai21  g564(.a(new_n411_), .b(new_n396_), .c(c), .O(new_n587_));
  gate1 g565(new_n587_, new_n586_, 1'b0, 1'b0, 1'b0, 1'b1, new_n588_);
  gate1 g566(n, new_n26_, 1'b0, 1'b0, 1'b0, d, new_n589_);
  gate1 g567(new_n589_, new_n63_, 1'b0, 1'b1, 1'b1, 1'b1, new_n590_);
  gate1 g568(new_n590_, new_n573_, 1'b0, 1'b0, 1'b0, 1'b1, new_n591_);
  gate1 g569(new_n591_, new_n588_, 1'b0, 1'b1, 1'b1, 1'b1, new_n592_);
  gate1 g570(new_n419_, new_n381_, 1'b0, 1'b0, 1'b0, 1'b1, new_n593_);
  oai21  g571(.a(new_n419_), .b(new_n381_), .c(c), .O(new_n594_));
  gate1 g572(new_n594_, new_n593_, 1'b0, 1'b0, 1'b0, 1'b1, new_n595_);
  gate1 g573(new_n595_, new_n541_, 1'b1, 1'b0, 1'b0, 1'b0, new_n596_);
  gate1 g574(new_n285_, new_n27_, d, 1'b1, 1'b1, 1'b1, new_n597_);
  gate1 g575(new_n597_, new_n596_, 1'b0, 1'b0, 1'b0, 1'b1, new_n598_);
  gate1 g576(n, d, 1'b1, 1'b1, 1'b1, 1'b0, new_n599_);
  gate1 g577(new_n595_, new_n552_, 1'b1, 1'b0, 1'b0, 1'b0, new_n600_);
  gate1 g578(new_n600_, new_n599_, 1'b0, 1'b0, 1'b0, new_n286_, new_n601_);
  gate1 g579(new_n558_, new_n416_, 1'b0, 1'b1, 1'b1, 1'b1, new_n602_);
  gate1 g580(new_n404_, new_n433_, 1'b0, 1'b0, 1'b0, new_n130_, new_n603_);
  gate1 g581(new_n558_, new_n603_, 1'b0, 1'b0, 1'b0, new_n262_, new_n604_);
  gate1 g582(new_n426_, new_n437_, 1'b0, 1'b0, 1'b0, 1'b1, new_n605_);
  gate1 g583(new_n541_, new_n605_, 1'b0, 1'b1, 1'b1, 1'b1, new_n606_);
  gate1 g584(new_n275_, new_n27_, 1'b0, 1'b1, 1'b1, 1'b1, new_n607_);
  gate1 g585(new_n607_, new_n541_, 1'b0, 1'b0, 1'b0, new_n605_, new_n608_);
  gate1 g586(new_n136_, new_n27_, l, 1'b1, 1'b1, 1'b1, new_n609_);
  gate1 g587(new_n441_, new_n109_, new_n27_, 1'b1, 1'b1, 1'b1, new_n610_);
  gate1 g588(new_n26_, d, 1'b0, 1'b1, 1'b1, 1'b1, new_n611_);
  gate1 g589(l, d, 1'b1, 1'b1, 1'b1, 1'b0, new_n612_);
  gate1 g590(new_n612_, new_n441_, 1'b0, 1'b0, 1'b0, new_n290_, new_n613_);
  gate1 g591(new_n296_, new_n26_, 1'b0, 1'b0, 1'b0, h, new_n614_);
  gate1 g592(new_n599_, new_n55_, 1'b0, 1'b0, 1'b0, new_n170_, new_n615_);
  gate1 g593(new_n615_, new_n614_, 1'b0, 1'b0, 1'b0, new_n613_, new_n616_);
  gate1 g594(new_n611_, ew_n610_), .c(new_n616_, 1'b0, 1'b1, new_n610_, 1'b1, new_n617_);
  gate1 g595(new_n447_, ew_n361_), .c(new_n358_, 1'b0, 1'b1, new_n361_, 1'b1, new_n618_);
  gate1 g596(new_n536_, new_n296_, 1'b0, 1'b0, 1'b0, l, new_n619_);
  gate1 g597(new_n619_, new_n618_, 1'b0, 1'b1, 1'b1, 1'b1, new_n620_);
  gate1 g598(new_n296_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n621_);
  gate1 g599(new_n621_, h, new_n529_, 1'b1, 1'b1, 1'b1, new_n622_);
  gate1 g600(new_n622_, ew_n618_), .c(new_n620_, 1'b0, 1'b1, new_n618_, 1'b1, new_n623_);
  gate1 g601(new_n530_, new_n295_, new_n27_, 1'b1, 1'b1, 1'b1, new_n624_);
  gate1 g602(new_n618_, new_n553_, new_n621_, 1'b1, 1'b1, 1'b1, new_n625_);
  gate1 g603(new_n624_, ew_n618_), .c(new_n625_, 1'b0, 1'b1, new_n618_, 1'b1, new_n626_);
  gate1 g604(new_n626_, new_n623_, 1'b0, 1'b0, 1'b0, new_n617_, new_n627_);
  gate1 g605(new_n609_, ew_n541_), .c(new_n627_, 1'b0, 1'b1, new_n541_, 1'b1, new_n628_);
  gate1 g606(new_n628_, new_n608_, 1'b0, 1'b0, 1'b0, 1'b1, new_n629_);
  gate1 g607(new_n606_, ew_n436_), .c(new_n629_, 1'b0, 1'b1, new_n436_, 1'b1, new_n630_);
  gate1 g608(new_n630_, new_n604_, 1'b0, 1'b0, 1'b0, 1'b1, new_n631_);
  gate1 g609(new_n631_, new_n602_, 1'b0, 1'b1, 1'b1, 1'b1, new_n632_);
  gate1 g610(new_n632_, new_n601_, 1'b0, 1'b0, 1'b0, new_n598_, new_n633_);
  gate1 g611(new_n194_, i, d, 1'b1, 1'b1, 1'b1, new_n634_);
  gate1 g612(new_n634_, new_n588_, 1'b0, 1'b0, 1'b0, new_n573_, new_n635_);
  gate1 g613(new_n590_, new_n588_, 1'b0, 1'b0, 1'b0, new_n558_, new_n636_);
  gate1 g614(new_n634_, new_n558_, 1'b1, 1'b1, 1'b1, 1'b0, new_n637_);
  gate1 g615(new_n637_, new_n587_, 1'b0, 1'b0, 1'b0, new_n586_, new_n638_);
  gate1 g616(new_n638_, new_n636_, 1'b0, 1'b0, 1'b0, new_n635_, new_n639_);
  gate1 g617(new_n639_, new_n633_, new_n592_, 1'b1, 1'b1, 1'b1, new_n640_);
  gate1 g618(new_n509_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n641_);
  gate1 g619(new_n561_, new_n560_, 1'b0, 1'b0, 1'b0, new_n573_, new_n642_);
  gate1 g620(new_n642_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n643_);
  gate1 g621(new_n562_, new_n560_, new_n573_, 1'b1, 1'b1, 1'b1, new_n644_);
  oai21  g622(.a(new_n644_), .b(new_n643_), .c(new_n641_), .O(new_n645_));
  gate1 g623(new_n645_, new_n640_, 1'b0, 1'b0, 1'b0, new_n585_, new_n646_);
  gate1 g624(new_n480_, new_n324_, 1'b0, 1'b0, 1'b0, new_n323_, new_n647_);
  gate1 g625(new_n647_, new_n646_, 1'b0, 1'b0, 1'b0, n, new_n648_);
  gate1 g626(new_n633_, new_n592_, 1'b0, 1'b1, 1'b1, 1'b1, new_n649_);
  gate1 g627(new_n639_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n650_);
  gate1 g628(new_n645_, new_n650_, 1'b0, 1'b0, 1'b0, new_n649_, new_n651_);
  gate1 g629(new_n651_, new_n584_, 1'b0, 1'b1, 1'b1, 1'b1, new_n652_);
  gate1 g630(new_n478_, new_n474_, new_n465_, 1'b1, 1'b1, 1'b1, new_n653_);
  gate1 g631(new_n653_, ew_n407_), .c(new_n481_, 1'b0, 1'b1, new_n407_, 1'b1, new_n654_);
  gate1 g632(new_n654_, new_n652_, 1'b0, 1'b0, 1'b0, n, new_n655_);
  gate1 g633(n, new_n510_, 1'b0, 1'b1, 1'b1, 1'b1, new_n656_);
  gate1 g634(new_n656_, new_n23_, 1'b0, 1'b0, 1'b0, new_n529_, new_n657_);
  gate1 g635(new_n27_, new_n23_, 1'b0, 1'b0, 1'b0, new_n510_, new_n658_);
  oai22  g636(.a(new_n658_), .b(new_n73_), .c(new_n657_), .d(new_n163_), .O(new_n659_));
  gate1 g637(new_n612_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n660_);
  gate1 g638(new_n656_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n661_);
  oai22  g639(.a(new_n658_), .b(new_n660_), .c(new_n661_), .d(new_n490_), .O(new_n662_));
  gate1 g640(new_n662_, new_n659_, 1'b0, 1'b1, 1'b1, 1'b1, new_n663_);
  gate1 g641(t, ew_n167_), .c(new_n178_, 1'b0, 1'b1, new_n167_, 1'b1, new_n664_);
  aoi22  g642(.a(new_n612_), .b(new_n169_), .c(new_n536_), .d(new_n335_), .O(new_n665_));
  gate1 g643(new_n665_, new_n664_, 1'b0, 1'b0, 1'b0, new_n663_, new_n666_);
  gate1 g644(new_n552_, ew_n183_), .c(new_n666_, 1'b0, 1'b1, new_n183_, 1'b1, new_n667_);
  gate1 g645(new_n36_, new_n510_, 1'b0, 1'b1, 1'b1, 1'b1, new_n668_);
  oai22  g646(.a(new_n668_), .b(new_n154_), .c(new_n550_), .d(new_n545_), .O(new_n669_));
  gate1 g647(new_n669_, new_n667_, 1'b0, 1'b0, 1'b0, 1'b1, new_n670_);
  gate1 g648(new_n570_, ew_n150_), .c(new_n670_, 1'b0, 1'b1, new_n150_, 1'b1, new_n671_);
  gate1 g649(new_n671_, new_n655_, 1'b0, 1'b0, 1'b0, new_n648_, r);
  gate1 g650(h, d, 1'b1, 1'b0, 1'b0, 1'b0, new_n673_);
  gate1 g651(new_n673_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, s);
  gate1 g652(new_n654_, new_n646_, 1'b0, 1'b0, 1'b0, n, new_n675_);
  gate1 g653(new_n173_, new_n27_, l, 1'b1, 1'b1, 1'b1, new_n676_);
  gate1 g654(new_n676_, i, 1'b1, 1'b1, 1'b1, 1'b0, new_n677_);
  gate1 g655(new_n677_, new_n580_, 1'b0, 1'b0, 1'b0, new_n541_, new_n678_);
  gate1 g656(new_n676_, new_n35_, 1'b0, 1'b0, 1'b0, 1'b1, new_n679_);
  gate1 g657(new_n679_, new_n573_, 1'b0, 1'b1, 1'b1, 1'b1, new_n680_);
  gate1 g658(new_n680_, new_n588_, 1'b0, 1'b0, 1'b0, 1'b1, new_n681_);
  gate1 g659(new_n676_, new_n35_, 1'b0, 1'b0, 1'b0, d, new_n682_);
  gate1 g660(new_n587_, ew_n586_), .c(new_n682_, 1'b0, 1'b1, new_n586_, 1'b1, new_n683_);
  gate1 g661(new_n560_, new_n558_, 1'b0, 1'b0, 1'b0, new_n137_, new_n684_);
  gate1 g662(new_n135_, new_n56_, new_n25_, 1'b1, 1'b1, 1'b1, new_n685_);
  gate1 g663(new_n685_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n686_);
  gate1 g664(new_n540_, ew_n525_), .c(new_n686_, 1'b0, 1'b1, new_n525_, 1'b1, new_n687_);
  gate1 g665(new_n606_, new_n272_, 1'b0, 1'b0, 1'b0, n, new_n688_);
  gate1 g666(new_n41_, new_n23_, i, 1'b1, 1'b1, 1'b1, new_n689_);
  gate1 g667(new_n689_, new_n606_, 1'b0, 1'b0, 1'b0, n, new_n690_);
  gate1 g668(new_n135_, new_n63_, 1'b0, 1'b1, 1'b1, 1'b1, new_n691_);
  gate1 g669(new_n691_, new_n541_, 1'b0, 1'b0, 1'b0, d, new_n692_);
  gate1 g670(new_n685_, new_n541_, 1'b0, 1'b0, 1'b0, d, new_n693_);
  gate1 g671(new_n618_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n694_);
  gate1 g672(new_n536_, new_n295_, new_n135_, 1'b1, 1'b1, 1'b1, new_n695_);
  gate1 g673(t, new_n456_, 1'b0, 1'b0, 1'b0, new_n134_, new_n696_);
  gate1 g674(new_n27_, new_n26_, d, 1'b1, 1'b1, 1'b1, new_n697_);
  gate1 g675(new_n697_, new_n442_, 1'b0, 1'b0, 1'b0, new_n110_, new_n698_);
  gate1 g676(new_n272_, n, 1'b0, 1'b0, 1'b0, new_n26_, new_n699_);
  gate1 g677(new_n699_, new_n698_, 1'b0, 1'b0, 1'b0, new_n696_, new_n700_);
  gate1 g678(new_n695_, ew_n694_), .c(new_n700_, 1'b0, 1'b1, new_n694_, 1'b1, new_n701_);
  gate1 g679(new_n701_, new_n693_, 1'b0, 1'b0, 1'b0, new_n692_, new_n702_);
  gate1 g680(new_n702_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n703_);
  gate1 g681(new_n703_, new_n690_, 1'b0, 1'b0, 1'b0, new_n688_, new_n704_);
  gate1 g682(new_n687_, ew_n595_), .c(new_n704_, 1'b0, 1'b1, new_n595_, 1'b1, new_n705_);
  gate1 g683(new_n685_, d, 1'b1, 1'b1, 1'b1, 1'b0, new_n706_);
  aoi22  g684(.a(new_n706_), .b(new_n595_), .c(new_n680_), .d(d), .O(new_n707_));
  gate1 g685(new_n707_, new_n705_, 1'b0, 1'b0, 1'b0, new_n684_, new_n708_);
  gate1 g686(new_n677_, new_n560_, 1'b0, 1'b0, 1'b0, new_n541_, new_n709_);
  gate1 g687(new_n603_, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, new_n710_);
  gate1 g688(new_n55_, new_n27_, l, 1'b1, 1'b1, 1'b1, new_n711_);
  gate1 g689(new_n711_, new_n573_, 1'b0, 1'b0, 1'b0, new_n710_, new_n712_);
  gate1 g690(new_n691_, new_n541_, 1'b1, 1'b1, 1'b1, 1'b0, new_n713_);
  gate1 g691(new_n135_, new_n63_, new_n529_, 1'b1, 1'b1, 1'b1, new_n714_);
  oai21  g692(.a(new_n714_), .b(new_n713_), .c(new_n595_), .O(new_n715_));
  gate1 g693(new_n715_, new_n712_, 1'b0, 1'b0, 1'b0, new_n709_, new_n716_);
  gate1 g694(new_n716_, new_n708_, new_n683_, 1'b1, 1'b1, 1'b1, new_n717_);
  gate1 g695(new_n717_, new_n681_, 1'b0, 1'b0, 1'b0, new_n678_, new_n718_);
  gate1 g696(new_n558_, new_n509_, 1'b0, 1'b0, 1'b0, new_n137_, new_n719_);
  gate1 g697(new_n677_, new_n580_, 1'b0, 1'b0, 1'b0, new_n560_, new_n720_);
  gate1 g698(new_n560_, new_n509_, 1'b0, 1'b0, 1'b0, new_n137_, new_n721_);
  gate1 g699(new_n721_, new_n720_, 1'b0, 1'b0, 1'b0, new_n719_, new_n722_);
  gate1 g700(new_n722_, new_n718_, 1'b0, 1'b1, 1'b1, 1'b1, new_n723_);
  gate1 g701(new_n723_, new_n675_, 1'b0, 1'b0, 1'b0, 1'b1, u);
  gate1 g702(new_n361_, new_n190_, new_n33_, 1'b1, 1'b1, 1'b1, new_n725_);
  gate1 g703(new_n673_, new_n371_, new_n362_, 1'b1, 1'b1, 1'b1, new_n726_);
  aoi22  g704(.a(new_n726_), .b(new_n297_), .c(new_n725_), .d(s), .O(new_n727_));
  gate1 g705(new_n190_, new_n33_, 1'b0, 1'b1, 1'b1, 1'b1, new_n728_);
  oai21  g706(.a(new_n728_), .b(new_n304_), .c(new_n726_), .O(new_n729_));
  gate1 g707(s, new_n197_, 1'b0, 1'b0, 1'b0, new_n32_, new_n730_);
  gate1 g708(new_n292_, new_n371_, 1'b0, 1'b0, 1'b0, new_n362_, new_n731_);
  gate1 g709(new_n292_, g, 1'b0, 1'b0, 1'b0, c, new_n732_);
  gate1 g710(new_n732_, ew_n731_), .c(new_n730_, 1'b0, 1'b1, new_n731_, 1'b1, new_n733_);
  gate1 g711(new_n360_, new_n334_, 1'b0, 1'b0, 1'b0, new_n49_, new_n734_);
  gate1 g712(new_n360_, new_n191_, 1'b0, 1'b0, 1'b0, new_n49_, new_n735_);
  gate1 g713(new_n735_, ew_n734_), .c(new_n673_, 1'b0, 1'b1, new_n734_, 1'b1, new_n736_);
  gate1 g714(new_n736_, new_n733_, 1'b0, 1'b1, 1'b1, 1'b1, new_n737_);
  gate1 g715(new_n737_, new_n729_, 1'b0, 1'b0, 1'b0, new_n727_, v);
endmodule


