// IWLS benchmark module "alu4_cl" printed on Wed May 29 16:26:22 2002
module test1(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n;
output
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v;
wire
  \[5] ,
  \[6] ,
  \[7] ,
  a1,
  a2,
  a3,
  a4,
  b1,
  b2,
  b3,
  b4,
  c1,
  c2,
  c3,
  c4,
  d1,
  d2,
  d3,
  d4,
  e1,
  e2,
  e3,
  e4,
  f1,
  f2,
  f3,
  f4,
  g1,
  g2,
  g3,
  g4,
  h1,
  h2,
  h3,
  h4,
  i1,
  i2,
  i3,
  i4,
  j1,
  j2,
  j3,
  j4,
  k1,
  k2,
  k3,
  k4,
  l1,
  l2,
  l3,
  l4,
  m0,
  m1,
  m2,
  m3,
  n0,
  n1,
  n2,
  n3,
  o0,
  o1,
  o2,
  o3,
  p0,
  p1,
  p2,
  p3,
  q0,
  q1,
  q2,
  q3,
  r0,
  r1,
  r2,
  r3,
  s0,
  s1,
  s2,
  s3,
  t0,
  t1,
  t2,
  t3,
  u0,
  u1,
  u2,
  u3,
  v0,
  v1,
  v2,
  v3,
  \[0] ,
  w0,
  w1,
  w2,
  w3,
  \[1] ,
  x0,
  x1,
  x2,
  x3,
  \[2] ,
  y0,
  y1,
  y2,
  y3,
  \[3] ,
  z0,
  z1,
  z2,
  z3,
  \[4] ;
assign
  \[5]  = h & d,
  \[6]  = (i1 & (h1 & (i & (s0 & (~l & n))))) | ((i1 & (z0 & (i & (s0 & (~l & n))))) | ((h1 & (c1 & (k & (~q0 & (l & n))))) | ((h1 & (z0 & (i & (s0 & (~l & n))))) | ((g1 & (d & (~i & (s0 & (~l & n))))) | ((g1 & (~i & (t0 & (s0 & (~l & n))))) | ((c1 & (d & (k & (~q0 & (l & n))))) | ((d & (~i & (t0 & (s0 & (~l & n))))) | ((h1 & (f1 & (c1 & (l & n)))) | ((f1 & (c1 & (d & (l & n)))) | ((e1 & (~d1 & (w0 & (l & n)))) | ((b1 & (k & (~q0 & (l & n)))) | ((a1 & (z0 & (x0 & (l & n)))) | ((a1 & (x0 & (t0 & (l & n)))) | ((z0 & (x0 & (t0 & (l & n)))) | ((~d & (y0 & (v0 & (l & n)))) | ((k & (r0 & (~l & (n0 & n)))) | ((u0 & (~t0 & (q0 & (~l & n)))) | ((f1 & (b1 & (l & n))) | ((\[5]  & (w0 & (l & n))) | ((~l & (o0 & n)) | ((p0 & (~m0 & n)) | (o0 & (n0 & n))))))))))))))))))))))),
  \[7]  = (~g & (y0 & (~f & (~e & \[4] )))) | ((d3 & (a2 & (~f & (~e & \[4] )))) | ((~z1 & (p2 & (k3 & \[4] ))) | ((~z1 & (k3 & (q2 & \[4] ))) | ((~z1 & (q2 & (j3 & \[4] ))) | ((p2 & (k3 & (a2 & \[4] ))) | ((k3 & (q2 & (a2 & \[4] ))) | (q2 & (j3 & (a2 & \[4] ))))))))),
  o = \[0] ,
  p = \[1] ,
  q = \[2] ,
  r = \[3] ,
  s = \[4] ,
  t = \[5] ,
  u = \[6] ,
  v = \[7] ,
  a1 = (w2 & u2) | ((w2 & v2) | (u2 & v2)),
  a2 = g & c,
  a3 = (~v2 & x3) | (v2 & ~x3),
  a4 = q3 & a,
  b1 = h1 & d,
  b2 = (o0 & l) | (q1 & j),
  b3 = (b & l3) | ((b & m2) | (l3 & m2)),
  b4 = u3 & n,
  c1 = (c & b3) | ((c & y1) | (b3 & y1)),
  c2 = (o0 & l) | (r0 & ~l),
  c3 = k & ~i,
  c4 = p1 & (j & n),
  d1 = ~h & ~d,
  d2 = u3 & ~j,
  d3 = ~b & ~a,
  d4 = (o1 & (~n & (l & ~j))) | ((r0 & (~u3 & n)) | (q0 & u3)),
  e1 = (z1 & t2) | a2,
  e2 = ~y1 & f3,
  e3 = ~q3 & ~r3,
  e4 = (l4 & (~n & v3)) | (n & (k & v3)),
  f1 = ~j & ~i,
  f2 = (~h1 & c1) | (h1 & ~c1),
  f3 = ~i3 & ~m2,
  f4 = (q0 & (l & ~k)) | (f1 & (l & ~k)),
  g1 = (c & x3) | ((c & v2) | (x3 & v2)),
  g2 = (~q0 & (k & l)) | (f1 & l),
  g3 = (~w3 & (i & (k & (i3 & (r2 & n))))) | ((w3 & (i & (k & (~i3 & (r2 & n))))) | ((~i & (~a & (k & (q3 & (r2 & n))))) | ((a & (l & (k & (~i3 & (~q0 & n))))) | ((~j & (a & (~i3 & (m1 & n)))) | ((j & (~l & (i3 & (m1 & n)))) | ((k1 & (~a & (l & (i3 & n)))) | ((~w3 & (x0 & (l & (q3 & n)))) | ((w3 & (x0 & (l & (~q3 & n)))) | ((~i & (a & (~q3 & (r2 & n)))) | ((n3 & (~k & (v3 & n))) | ((m3 & (~k & (v3 & n))) | ((v0 & (~a & (l & n))) | ((e & (x2 & (r2 & n))) | ((a & (~l & (m1 & n))) | ((~q3 & (q0 & (u3 & n))) | (~i3 & (b2 & n))))))))))))))))),
  g4 = (~g & c) | ((~g & ~j4) | (c & ~j4)),
  h1 = (j & (u3 & (g4 & (~d & (~i & (n & h)))))) | ((j & (g4 & (d & (~i & (n & ~h))))) | ((~l & (~k & (~d & (~i & ~n)))) | ((~j & (~k & (~d & (~i & ~n)))) | ((j & (~g4 & (~i & (n & d1)))) | ((u3 & (~g4 & (~i & (n & \[5] )))) | ((s0 & (x1 & (~i & n))) | ((f4 & (n & \[5] )) | ((d2 & (~i & \[5] )) | ((d2 & (n & \[5] )) | ((~h & d4) | (e4 & ~d1))))))))))),
  h2 = (~h1 & z0) | (h1 & ~z0),
  h3 = l & a,
  h4 = (d2 & n) | k4,
  i1 = (z2 & u2) | ((z2 & y1) | (u2 & y1)),
  i2 = (f1 & ~k) | g2,
  i3 = (n3 & (u3 & (n & r0))) | ((m3 & (n & r0)) | ((~e & d4) | ((~a & i4) | ((k3 & k4) | (e4 & ~j3))))),
  i4 = (~l & (~n & m1)) | (~j & (~n & m1)),
  j1 = (q0 & (l4 & n)) | (s0 & (p1 & ~n)),
  j2 = ~q0 & l4,
  j3 = ~e & ~a,
  j4 = (n3 & ~n2) | o2,
  k1 = f1 | k,
  k2 = ~g3 | m,
  k3 = e & a,
  k4 = (q1 & ~j) | (f4 & n),
  l1 = l & d,
  l2 = (~s3 & (~p3 & (o1 & (m2 & (r2 & n))))) | ((~s3 & (p3 & (o1 & (~m2 & (r2 & n))))) | ((s3 & (~p3 & (o1 & (~m2 & (r2 & n))))) | ((s3 & (p3 & (o1 & (m2 & (r2 & n))))) | ((p2 & (k3 & (l & (w0 & n)))) | ((~k3 & (~f & (b & (w0 & n)))) | ((i2 & (b & (~l3 & (~m2 & n)))) | ((i2 & (b & (l3 & (m2 & n)))) | ((~t3 & (~s3 & (r3 & (s2 & n)))) | ((~t3 & (s3 & (~r3 & (s2 & n)))) | ((t3 & (~s3 & (~r3 & (s2 & n)))) | ((t3 & (s3 & (r3 & (s2 & n)))) | ((r3 & (q3 & (~l & (v0 & n)))) | ((~i & (~o3 & (b & (r2 & n)))) | ((c3 & (o3 & (~b & (r2 & n)))) | ((~b & (~l3 & (m2 & (g2 & n)))) | ((~b & (l3 & (~m2 & (g2 & n)))) | ((q2 & (k3 & (w0 & n))) | ((o2 & (~k3 & (w0 & n))) | ((i3 & (c2 & (m2 & n))) | ((x0 & (~l & (m2 & n))) | ((h3 & (b & (v0 & n))) | ((e3 & (~l & (v0 & n))) | ((l & (d3 & (v0 & n))) | ((f & (x2 & (r2 & n))) | ((j2 & (b & n)) | (f3 & (b2 & n))))))))))))))))))))))))))),
  l3 = i3 & a,
  l4 = ~l & ~k,
  m0 = ~w1 | v1,
  m1 = ~k & ~i,
  m2 = (o2 & (j & (~n3 & (u3 & (~i & n))))) | ((n2 & (j & (~n3 & (~i & n)))) | ((j & (n3 & (~i & (n & p2)))) | ((n3 & (u3 & (~i & (n & q2)))) | ((h3 & (s0 & (~i & n))) | ((~f & d4) | ((~b & i4) | ((q2 & h4) | (e4 & ~p2)))))))),
  m3 = ~e & a,
  n0 = e2 & ~h1,
  n1 = c3 | l,
  n2 = ~f & b,
  n3 = e & ~a,
  o0 = q0 & ~k,
  o1 = k & i,
  o2 = f & ~b,
  o3 = (~a4 & r3) | (a4 & ~r3),
  p0 = (f1 & (~g1 & (~t0 & (~l & (d & n))))) | ((f1 & (g1 & (t0 & (~l & (d & n))))) | ((~g1 & (t0 & (~i & (~d & (d2 & n))))) | ((g1 & (~t0 & (~i & (~d & (d2 & n))))) | ((~a1 & (~t0 & (z0 & (l & (x0 & n))))) | ((~a1 & (t0 & (~z0 & (l & (x0 & n))))) | ((a1 & (~t0 & (~z0 & (l & (x0 & n))))) | ((a1 & (t0 & (z0 & (l & (x0 & n))))) | ((d1 & (e1 & (l & (w0 & n)))) | ((~i1 & (h2 & (i & (d2 & n)))) | ((i1 & (~h2 & (i & (d2 & n)))) | ((~u0 & (t0 & (~l & (v0 & n)))) | ((u0 & (~t0 & (~l & (v0 & n)))) | ((~h & (~e1 & (d & (w0 & n)))) | ((h & (~e1 & (~d & (w0 & n)))) | ((l & (~d & (y0 & (v0 & n)))) | ((\[5]  & (e1 & (w0 & n))) | ((i2 & (~f2 & (d & n))) | ((h & (~l & (w0 & n))) | ((g2 & (f2 & (~d & n))) | ((~l & (h1 & (x0 & n))) | ((~y0 & (l1 & (v0 & n))) | ((~e2 & (h1 & (c2 & n))) | ((j2 & (d & n)) | (n0 & (b2 & n))))))))))))))))))))))))),
  p1 = l & ~i,
  p2 = ~f & ~b,
  p3 = i3 & w3,
  q0 = j & i,
  q1 = u3 & ~i,
  q2 = f & b,
  q3 = (v3 & (k3 & b4)) | ((q0 & (l3 & b4)) | ((f1 & (~i3 & b4)) | ((a & c4) | (i3 & c4)))),
  r0 = j & ~i,
  r1 = (l & k) | m1,
  r2 = ~l & ~j,
  r3 = (~j & (f & (i & (b & b4)))) | ((j & (i & (b & (m2 & b4)))) | ((~m2 & (f1 & b4)) | ((b & c4) | (m2 & c4)))),
  s0 = k & ~j,
  s1 = (l4 & i) | c3,
  s2 = p1 & (j & ~k),
  s3 = (q2 & y3) | (z3 & ~r3),
  t0 = (v3 & (\[5]  & b4)) | ((q0 & (b1 & b4)) | ((f1 & (~h1 & b4)) | ((d & c4) | (h1 & c4)))),
  t1 = x2 & l,
  t2 = (~p2 & k3) | q2,
  t3 = q3 & w3,
  u0 = ~v2 & e3,
  u1 = u3 & i,
  u2 = (a2 & y3) | (z3 & ~v2),
  u3 = ~l & k,
  v0 = q0 & k,
  v1 = ~l2 | k2,
  v2 = (~j & (g & (i & (c & b4)))) | ((j & (i & (c & (y1 & b4)))) | ((~y1 & (f1 & b4)) | ((c & c4) | (y1 & c4)))),
  v3 = ~j & i,
  \[0]  = (n3 & (t1 & (~j & ~n))) | ((m3 & (l & (~j & ~n))) | ((u1 & (~j & (~e & ~n))) | ((r1 & (~j & (i3 & ~n))) | ((s1 & (~j & (~i3 & ~n))) | ((l3 & (o1 & (j & ~n))) | ((k3 & (n1 & (j & ~n))) | ((q1 & (j3 & (j & ~n))) | ((p1 & (j & (e & ~n))) | ((e & (i3 & (m1 & ~n))) | ((h3 & (k1 & ~n)) | ((~m & (~g3 & n)) | ((m & (g3 & n)) | j1)))))))))))),
  w0 = x2 & ~j,
  w1 = (~z1 & (l & (t2 & (w0 & n)))) | ((~e3 & (~l & (v2 & (v0 & n)))) | ((c3 & (a3 & (~c & (r2 & n)))) | ((g2 & (~b3 & (~c & (y1 & n)))) | ((g2 & (b3 & (~c & (~y1 & n)))) | ((~b3 & (i2 & (c & (~y1 & n)))) | ((b3 & (i2 & (c & (y1 & n)))) | ((~i & (~a3 & (c & (r2 & n)))) | ((~z2 & (~y2 & (o1 & (r2 & n)))) | ((z2 & (y2 & (o1 & (r2 & n)))) | ((~g & (c & (~t2 & (w0 & n)))) | ((g & (~c & (~t2 & (w0 & n)))) | ((~w2 & (~v2 & (u2 & (s2 & n)))) | ((~w2 & (v2 & (~u2 & (s2 & n)))) | ((w2 & (~v2 & (~u2 & (s2 & n)))) | ((w2 & (v2 & (u2 & (s2 & n)))) | ((a2 & (t2 & (w0 & n))) | ((~f3 & (c2 & (y1 & n))) | ((x0 & (~l & (y1 & n))) | ((u0 & (~l & (v0 & n))) | ((l & (y0 & (v0 & n))) | ((~d3 & (x1 & (v0 & n))) | ((g & (x2 & (r2 & n))) | ((j2 & (c & n)) | (e2 & (b2 & n))))))))))))))))))))))))),
  w2 = (t3 & s3) | ((t3 & r3) | (s3 & r3)),
  w3 = (k3 & y3) | (z3 & ~q3),
  \[1]  = (o1 & (j & (b & (m2 & ~n)))) | ((q2 & (n1 & (j & ~n))) | ((p2 & (q1 & (j & ~n))) | ((p1 & (j & (f & ~n))) | ((o2 & (t1 & (~j & ~n))) | ((n2 & (l & (~j & ~n))) | ((u1 & (~j & (~f & ~n))) | ((r1 & (~j & (m2 & ~n))) | ((s1 & (~j & (~m2 & ~n))) | ((l & (b & (k1 & ~n))) | ((f & (m2 & (m1 & ~n))) | ((~l2 & (~k2 & n)) | ((l2 & (k2 & n)) | j1)))))))))))),
  x0 = m1 & j,
  x1 = l & c,
  x2 = ~k & i,
  x3 = (b & a4) | ((b & r3) | (a4 & r3)),
  \[2]  = (t1 & (~c & (~j & (g & ~n)))) | ((c & (o1 & (j & (y1 & ~n)))) | ((u1 & (~j & (~g & ~n))) | ((s1 & (~j & (~y1 & ~n))) | ((r1 & (~j & (y1 & ~n))) | ((q1 & (~z1 & (j & ~n))) | ((p1 & (j & (g & ~n))) | ((a2 & (n1 & (j & ~n))) | ((~j & (~g & (x1 & ~n))) | ((g & (y1 & (m1 & ~n))) | ((x1 & (k1 & ~n)) | ((~w1 & (~v1 & n)) | ((w1 & (v1 & n)) | j1)))))))))))),
  y0 = d3 & ~c,
  y1 = (j & (~j4 & (u3 & (~i & (n & (g & ~c)))))) | ((j & (~j4 & (~i & (n & (~g & c))))) | ((j & (j4 & (~i & (n & (~g & ~c))))) | ((j4 & (u3 & (~i & (n & (g & c))))) | ((l & (b & (s0 & (~i & n)))) | ((~g & d4) | ((~c & i4) | ((e4 & z1) | (a2 & h4)))))))),
  y2 = (~y1 & ~u2) | (y1 & u2),
  y3 = c4 & ~k,
  \[3]  = (~d & (t1 & (~j & (h & ~n)))) | ((u1 & (~j & (~h & ~n))) | ((s1 & (~j & (~h1 & ~n))) | ((r1 & (~j & (h1 & ~n))) | ((\[5]  & (n1 & (j & ~n))) | ((d1 & (q1 & (j & ~n))) | ((b1 & (o1 & (j & ~n))) | ((p1 & (j & (h & ~n))) | ((~j & (~h & (l1 & ~n))) | ((h & (h1 & (m1 & ~n))) | ((l1 & (k1 & ~n)) | ((~p0 & (~m0 & n)) | ((p0 & (m0 & n)) | j1)))))))))))),
  z0 = (\[5]  & y3) | (z3 & ~t0),
  z1 = g | c,
  z2 = (p3 & s3) | ((p3 & m2) | (s3 & m2)),
  z3 = u1 & (n & ~j),
  \[4]  = d1 | \[5] ;
endmodule

